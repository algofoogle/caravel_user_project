VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_example
  CLASS BLOCK ;
  FOREIGN user_proj_example ;
  ORIGIN 0.000 0.000 ;
  SIZE 2700.000 BY 1500.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 31.320 2700.000 31.920 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1010.520 2700.000 1011.120 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1108.440 2700.000 1109.040 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1206.360 2700.000 1206.960 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1304.280 2700.000 1304.880 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1402.200 2700.000 1402.800 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2647.390 1496.000 2647.670 1500.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2347.930 1496.000 2348.210 1500.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2048.470 1496.000 2048.750 1500.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1749.010 1496.000 1749.290 1500.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1449.550 1496.000 1449.830 1500.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 129.240 2700.000 129.840 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1150.090 1496.000 1150.370 1500.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 850.630 1496.000 850.910 1500.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.170 1496.000 551.450 1500.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.710 1496.000 251.990 1500.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1474.280 4.000 1474.880 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1368.200 4.000 1368.800 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1262.120 4.000 1262.720 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1156.040 4.000 1156.640 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1049.960 4.000 1050.560 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 943.880 4.000 944.480 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 227.160 2700.000 227.760 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 837.800 4.000 838.400 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 731.720 4.000 732.320 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 625.640 4.000 626.240 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 519.560 4.000 520.160 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 413.480 4.000 414.080 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 307.400 4.000 308.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 201.320 4.000 201.920 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 325.080 2700.000 325.680 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 423.000 2700.000 423.600 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2696.000 520.920 2700.000 521.520 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2696.000 618.840 2700.000 619.440 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2696.000 716.760 2700.000 717.360 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2696.000 814.680 2700.000 815.280 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 2696.000 912.600 2700.000 913.200 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 96.600 2700.000 97.200 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1075.800 2700.000 1076.400 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1173.720 2700.000 1174.320 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1271.640 2700.000 1272.240 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1369.560 2700.000 1370.160 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1467.480 2700.000 1468.080 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2447.750 1496.000 2448.030 1500.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2148.290 1496.000 2148.570 1500.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1848.830 1496.000 1849.110 1500.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1549.370 1496.000 1549.650 1500.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1249.910 1496.000 1250.190 1500.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 194.520 2700.000 195.120 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 950.450 1496.000 950.730 1500.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.990 1496.000 651.270 1500.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.530 1496.000 351.810 1500.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.070 1496.000 52.350 1500.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1403.560 4.000 1404.160 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1297.480 4.000 1298.080 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1191.400 4.000 1192.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1085.320 4.000 1085.920 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 979.240 4.000 979.840 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 873.160 4.000 873.760 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 292.440 2700.000 293.040 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 767.080 4.000 767.680 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 661.000 4.000 661.600 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 554.920 4.000 555.520 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.840 4.000 449.440 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.760 4.000 343.360 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.680 4.000 237.280 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 4.000 131.200 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 4.000 25.120 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 390.360 2700.000 390.960 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 488.280 2700.000 488.880 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2696.000 586.200 2700.000 586.800 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2696.000 684.120 2700.000 684.720 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2696.000 782.040 2700.000 782.640 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2696.000 879.960 2700.000 880.560 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2696.000 977.880 2700.000 978.480 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2696.000 63.960 2700.000 64.560 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1043.160 2700.000 1043.760 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1141.080 2700.000 1141.680 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1239.000 2700.000 1239.600 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1336.920 2700.000 1337.520 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1434.840 2700.000 1435.440 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2547.570 1496.000 2547.850 1500.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2248.110 1496.000 2248.390 1500.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1948.650 1496.000 1948.930 1500.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1649.190 1496.000 1649.470 1500.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1349.730 1496.000 1350.010 1500.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2696.000 161.880 2700.000 162.480 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1050.270 1496.000 1050.550 1500.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 750.810 1496.000 751.090 1500.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 451.350 1496.000 451.630 1500.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 151.890 1496.000 152.170 1500.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1438.920 4.000 1439.520 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1332.840 4.000 1333.440 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1226.760 4.000 1227.360 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1120.680 4.000 1121.280 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1014.600 4.000 1015.200 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 908.520 4.000 909.120 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2696.000 259.800 2700.000 260.400 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 802.440 4.000 803.040 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 696.360 4.000 696.960 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 590.280 4.000 590.880 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 484.200 4.000 484.800 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.120 4.000 378.720 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 4.000 166.560 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 4.000 60.480 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2696.000 357.720 2700.000 358.320 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2696.000 455.640 2700.000 456.240 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2696.000 553.560 2700.000 554.160 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2696.000 651.480 2700.000 652.080 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2696.000 749.400 2700.000 750.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2696.000 847.320 2700.000 847.920 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2696.000 945.240 2700.000 945.840 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2581.610 0.000 2581.890 4.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2586.670 0.000 2586.950 4.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2591.730 0.000 2592.010 4.000 ;
    END
  END irq[2]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 638.570 0.000 638.850 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2156.570 0.000 2156.850 4.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2171.750 0.000 2172.030 4.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2186.930 0.000 2187.210 4.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2202.110 0.000 2202.390 4.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2217.290 0.000 2217.570 4.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2232.470 0.000 2232.750 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2247.650 0.000 2247.930 4.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2262.830 0.000 2263.110 4.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2278.010 0.000 2278.290 4.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2293.190 0.000 2293.470 4.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 790.370 0.000 790.650 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2308.370 0.000 2308.650 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2323.550 0.000 2323.830 4.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2338.730 0.000 2339.010 4.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2353.910 0.000 2354.190 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2369.090 0.000 2369.370 4.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2384.270 0.000 2384.550 4.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2399.450 0.000 2399.730 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2414.630 0.000 2414.910 4.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2429.810 0.000 2430.090 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2444.990 0.000 2445.270 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.550 0.000 805.830 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2460.170 0.000 2460.450 4.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2475.350 0.000 2475.630 4.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2490.530 0.000 2490.810 4.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2505.710 0.000 2505.990 4.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2520.890 0.000 2521.170 4.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2536.070 0.000 2536.350 4.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2551.250 0.000 2551.530 4.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2566.430 0.000 2566.710 4.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 820.730 0.000 821.010 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 835.910 0.000 836.190 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.090 0.000 851.370 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 866.270 0.000 866.550 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 881.450 0.000 881.730 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 896.630 0.000 896.910 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.810 0.000 912.090 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 926.990 0.000 927.270 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.750 0.000 654.030 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.170 0.000 942.450 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 957.350 0.000 957.630 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.530 0.000 972.810 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 987.710 0.000 987.990 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1002.890 0.000 1003.170 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1018.070 0.000 1018.350 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1033.250 0.000 1033.530 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1048.430 0.000 1048.710 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1063.610 0.000 1063.890 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1078.790 0.000 1079.070 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.930 0.000 669.210 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1093.970 0.000 1094.250 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1109.150 0.000 1109.430 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1124.330 0.000 1124.610 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1139.510 0.000 1139.790 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1154.690 0.000 1154.970 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1169.870 0.000 1170.150 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1185.050 0.000 1185.330 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1200.230 0.000 1200.510 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1215.410 0.000 1215.690 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1230.590 0.000 1230.870 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 684.110 0.000 684.390 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1245.770 0.000 1246.050 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1260.950 0.000 1261.230 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1276.130 0.000 1276.410 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.310 0.000 1291.590 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1306.490 0.000 1306.770 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1321.670 0.000 1321.950 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1336.850 0.000 1337.130 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1352.030 0.000 1352.310 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1367.210 0.000 1367.490 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1382.390 0.000 1382.670 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.290 0.000 699.570 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1397.570 0.000 1397.850 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1412.750 0.000 1413.030 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1427.930 0.000 1428.210 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1443.110 0.000 1443.390 4.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1458.290 0.000 1458.570 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1473.470 0.000 1473.750 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1488.650 0.000 1488.930 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1503.830 0.000 1504.110 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1519.010 0.000 1519.290 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1534.190 0.000 1534.470 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.470 0.000 714.750 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1549.370 0.000 1549.650 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1564.550 0.000 1564.830 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1579.730 0.000 1580.010 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1594.910 0.000 1595.190 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1610.090 0.000 1610.370 4.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1625.270 0.000 1625.550 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1640.450 0.000 1640.730 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1655.630 0.000 1655.910 4.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1670.810 0.000 1671.090 4.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1685.990 0.000 1686.270 4.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.650 0.000 729.930 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1701.170 0.000 1701.450 4.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1716.350 0.000 1716.630 4.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1731.530 0.000 1731.810 4.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1746.710 0.000 1746.990 4.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1761.890 0.000 1762.170 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1777.070 0.000 1777.350 4.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1792.250 0.000 1792.530 4.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1807.430 0.000 1807.710 4.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1822.610 0.000 1822.890 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1837.790 0.000 1838.070 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 744.830 0.000 745.110 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1852.970 0.000 1853.250 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1868.150 0.000 1868.430 4.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 1883.330 0.000 1883.610 4.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1898.510 0.000 1898.790 4.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1913.690 0.000 1913.970 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1928.870 0.000 1929.150 4.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1944.050 0.000 1944.330 4.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1959.230 0.000 1959.510 4.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1974.410 0.000 1974.690 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1989.590 0.000 1989.870 4.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.010 0.000 760.290 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2004.770 0.000 2005.050 4.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2019.950 0.000 2020.230 4.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2035.130 0.000 2035.410 4.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2050.310 0.000 2050.590 4.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2065.490 0.000 2065.770 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2080.670 0.000 2080.950 4.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2095.850 0.000 2096.130 4.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2111.030 0.000 2111.310 4.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2126.210 0.000 2126.490 4.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2141.390 0.000 2141.670 4.000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.190 0.000 775.470 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 643.630 0.000 643.910 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2161.630 0.000 2161.910 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2176.810 0.000 2177.090 4.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2191.990 0.000 2192.270 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2207.170 0.000 2207.450 4.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2222.350 0.000 2222.630 4.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2237.530 0.000 2237.810 4.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2252.710 0.000 2252.990 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2267.890 0.000 2268.170 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2283.070 0.000 2283.350 4.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2298.250 0.000 2298.530 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 795.430 0.000 795.710 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2313.430 0.000 2313.710 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2328.610 0.000 2328.890 4.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2343.790 0.000 2344.070 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2358.970 0.000 2359.250 4.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2374.150 0.000 2374.430 4.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2389.330 0.000 2389.610 4.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2404.510 0.000 2404.790 4.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2419.690 0.000 2419.970 4.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2434.870 0.000 2435.150 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2450.050 0.000 2450.330 4.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 810.610 0.000 810.890 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2465.230 0.000 2465.510 4.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2480.410 0.000 2480.690 4.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2495.590 0.000 2495.870 4.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2510.770 0.000 2511.050 4.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2525.950 0.000 2526.230 4.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2541.130 0.000 2541.410 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2556.310 0.000 2556.590 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2571.490 0.000 2571.770 4.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 825.790 0.000 826.070 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 840.970 0.000 841.250 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 856.150 0.000 856.430 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 871.330 0.000 871.610 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 886.510 0.000 886.790 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.690 0.000 901.970 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 916.870 0.000 917.150 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.050 0.000 932.330 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 658.810 0.000 659.090 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 947.230 0.000 947.510 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 962.410 0.000 962.690 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 977.590 0.000 977.870 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 992.770 0.000 993.050 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.950 0.000 1008.230 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1023.130 0.000 1023.410 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1038.310 0.000 1038.590 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1053.490 0.000 1053.770 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1068.670 0.000 1068.950 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1083.850 0.000 1084.130 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 673.990 0.000 674.270 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1099.030 0.000 1099.310 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1114.210 0.000 1114.490 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1129.390 0.000 1129.670 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1144.570 0.000 1144.850 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1159.750 0.000 1160.030 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1174.930 0.000 1175.210 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1190.110 0.000 1190.390 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1205.290 0.000 1205.570 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1220.470 0.000 1220.750 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1235.650 0.000 1235.930 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 689.170 0.000 689.450 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1250.830 0.000 1251.110 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1266.010 0.000 1266.290 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1281.190 0.000 1281.470 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1296.370 0.000 1296.650 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1311.550 0.000 1311.830 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1326.730 0.000 1327.010 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1341.910 0.000 1342.190 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1357.090 0.000 1357.370 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1372.270 0.000 1372.550 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1387.450 0.000 1387.730 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 704.350 0.000 704.630 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1402.630 0.000 1402.910 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1417.810 0.000 1418.090 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1432.990 0.000 1433.270 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1448.170 0.000 1448.450 4.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1463.350 0.000 1463.630 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1478.530 0.000 1478.810 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1493.710 0.000 1493.990 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1508.890 0.000 1509.170 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1524.070 0.000 1524.350 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1539.250 0.000 1539.530 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 719.530 0.000 719.810 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1554.430 0.000 1554.710 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1569.610 0.000 1569.890 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1584.790 0.000 1585.070 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1599.970 0.000 1600.250 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1615.150 0.000 1615.430 4.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1630.330 0.000 1630.610 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1645.510 0.000 1645.790 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1660.690 0.000 1660.970 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1675.870 0.000 1676.150 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1691.050 0.000 1691.330 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 734.710 0.000 734.990 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1706.230 0.000 1706.510 4.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1721.410 0.000 1721.690 4.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1736.590 0.000 1736.870 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1751.770 0.000 1752.050 4.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1766.950 0.000 1767.230 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1782.130 0.000 1782.410 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1797.310 0.000 1797.590 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1812.490 0.000 1812.770 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1827.670 0.000 1827.950 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1842.850 0.000 1843.130 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 749.890 0.000 750.170 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1858.030 0.000 1858.310 4.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1873.210 0.000 1873.490 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1888.390 0.000 1888.670 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1903.570 0.000 1903.850 4.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1918.750 0.000 1919.030 4.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1933.930 0.000 1934.210 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1949.110 0.000 1949.390 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1964.290 0.000 1964.570 4.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1979.470 0.000 1979.750 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1994.650 0.000 1994.930 4.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 765.070 0.000 765.350 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2009.830 0.000 2010.110 4.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2025.010 0.000 2025.290 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2040.190 0.000 2040.470 4.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2055.370 0.000 2055.650 4.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2070.550 0.000 2070.830 4.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2085.730 0.000 2086.010 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2100.910 0.000 2101.190 4.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2116.090 0.000 2116.370 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2131.270 0.000 2131.550 4.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2146.450 0.000 2146.730 4.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 780.250 0.000 780.530 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 648.690 0.000 648.970 4.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2166.690 0.000 2166.970 4.000 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2181.870 0.000 2182.150 4.000 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2197.050 0.000 2197.330 4.000 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2212.230 0.000 2212.510 4.000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2227.410 0.000 2227.690 4.000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2242.590 0.000 2242.870 4.000 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2257.770 0.000 2258.050 4.000 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2272.950 0.000 2273.230 4.000 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2288.130 0.000 2288.410 4.000 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2303.310 0.000 2303.590 4.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.490 0.000 800.770 4.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2318.490 0.000 2318.770 4.000 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2333.670 0.000 2333.950 4.000 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2348.850 0.000 2349.130 4.000 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2364.030 0.000 2364.310 4.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2379.210 0.000 2379.490 4.000 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2394.390 0.000 2394.670 4.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2409.570 0.000 2409.850 4.000 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2424.750 0.000 2425.030 4.000 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2439.930 0.000 2440.210 4.000 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2455.110 0.000 2455.390 4.000 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 815.670 0.000 815.950 4.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2470.290 0.000 2470.570 4.000 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2485.470 0.000 2485.750 4.000 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2500.650 0.000 2500.930 4.000 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2515.830 0.000 2516.110 4.000 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2531.010 0.000 2531.290 4.000 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2546.190 0.000 2546.470 4.000 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2561.370 0.000 2561.650 4.000 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2576.550 0.000 2576.830 4.000 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.850 0.000 831.130 4.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.030 0.000 846.310 4.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 861.210 0.000 861.490 4.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 876.390 0.000 876.670 4.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 891.570 0.000 891.850 4.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 906.750 0.000 907.030 4.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.930 0.000 922.210 4.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 937.110 0.000 937.390 4.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.870 0.000 664.150 4.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 952.290 0.000 952.570 4.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 967.470 0.000 967.750 4.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 982.650 0.000 982.930 4.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 997.830 0.000 998.110 4.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.010 0.000 1013.290 4.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1028.190 0.000 1028.470 4.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1043.370 0.000 1043.650 4.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1058.550 0.000 1058.830 4.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1073.730 0.000 1074.010 4.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1088.910 0.000 1089.190 4.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.050 0.000 679.330 4.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1104.090 0.000 1104.370 4.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1119.270 0.000 1119.550 4.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1134.450 0.000 1134.730 4.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1149.630 0.000 1149.910 4.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1164.810 0.000 1165.090 4.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1179.990 0.000 1180.270 4.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1195.170 0.000 1195.450 4.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1210.350 0.000 1210.630 4.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1225.530 0.000 1225.810 4.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1240.710 0.000 1240.990 4.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.230 0.000 694.510 4.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1255.890 0.000 1256.170 4.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1271.070 0.000 1271.350 4.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1286.250 0.000 1286.530 4.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1301.430 0.000 1301.710 4.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1316.610 0.000 1316.890 4.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1331.790 0.000 1332.070 4.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1346.970 0.000 1347.250 4.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1362.150 0.000 1362.430 4.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1377.330 0.000 1377.610 4.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1392.510 0.000 1392.790 4.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 709.410 0.000 709.690 4.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1407.690 0.000 1407.970 4.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1422.870 0.000 1423.150 4.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1438.050 0.000 1438.330 4.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1453.230 0.000 1453.510 4.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1468.410 0.000 1468.690 4.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1483.590 0.000 1483.870 4.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1498.770 0.000 1499.050 4.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1513.950 0.000 1514.230 4.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1529.130 0.000 1529.410 4.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1544.310 0.000 1544.590 4.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.590 0.000 724.870 4.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1559.490 0.000 1559.770 4.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1574.670 0.000 1574.950 4.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1589.850 0.000 1590.130 4.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1605.030 0.000 1605.310 4.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1620.210 0.000 1620.490 4.000 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1635.390 0.000 1635.670 4.000 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1650.570 0.000 1650.850 4.000 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1665.750 0.000 1666.030 4.000 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1680.930 0.000 1681.210 4.000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1696.110 0.000 1696.390 4.000 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 739.770 0.000 740.050 4.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1711.290 0.000 1711.570 4.000 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1726.470 0.000 1726.750 4.000 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1741.650 0.000 1741.930 4.000 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1756.830 0.000 1757.110 4.000 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1772.010 0.000 1772.290 4.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1787.190 0.000 1787.470 4.000 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1802.370 0.000 1802.650 4.000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1817.550 0.000 1817.830 4.000 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1832.730 0.000 1833.010 4.000 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1847.910 0.000 1848.190 4.000 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.950 0.000 755.230 4.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1863.090 0.000 1863.370 4.000 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1878.270 0.000 1878.550 4.000 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1893.450 0.000 1893.730 4.000 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1908.630 0.000 1908.910 4.000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1923.810 0.000 1924.090 4.000 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1938.990 0.000 1939.270 4.000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1954.170 0.000 1954.450 4.000 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1969.350 0.000 1969.630 4.000 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1984.530 0.000 1984.810 4.000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1999.710 0.000 1999.990 4.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.130 0.000 770.410 4.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2014.890 0.000 2015.170 4.000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2030.070 0.000 2030.350 4.000 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2045.250 0.000 2045.530 4.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2060.430 0.000 2060.710 4.000 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2075.610 0.000 2075.890 4.000 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2090.790 0.000 2091.070 4.000 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2105.970 0.000 2106.250 4.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2121.150 0.000 2121.430 4.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2136.330 0.000 2136.610 4.000 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2151.510 0.000 2151.790 4.000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.310 0.000 785.590 4.000 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2596.790 0.000 2597.070 4.000 ;
    END
  END user_clock2
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.640 10.640 1712.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.240 10.640 1865.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2017.840 10.640 2019.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2171.440 10.640 2173.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2325.040 10.640 2326.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2478.640 10.640 2480.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2632.240 10.640 2633.840 1488.080 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1787.440 10.640 1789.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1941.040 10.640 1942.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2094.640 10.640 2096.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2248.240 10.640 2249.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2401.840 10.640 2403.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2555.440 10.640 2557.040 1488.080 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 107.270 0.000 107.550 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 0.000 132.850 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.610 0.000 304.890 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.790 0.000 320.070 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 0.000 335.250 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.150 0.000 350.430 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.330 0.000 365.610 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.510 0.000 380.790 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.690 0.000 395.970 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.870 0.000 411.150 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.050 0.000 426.330 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.230 0.000 441.510 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.810 0.000 153.090 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.410 0.000 456.690 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.590 0.000 471.870 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.770 0.000 487.050 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.950 0.000 502.230 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.130 0.000 517.410 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.310 0.000 532.590 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 0.000 547.770 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.670 0.000 562.950 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.850 0.000 578.130 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.030 0.000 593.310 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.050 0.000 173.330 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.210 0.000 608.490 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.390 0.000 623.670 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.530 0.000 213.810 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.890 0.000 244.170 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.070 0.000 259.350 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.250 0.000 274.530 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.430 0.000 289.710 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 117.390 0.000 117.670 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 137.630 0.000 137.910 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 309.670 0.000 309.950 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 324.850 0.000 325.130 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 340.030 0.000 340.310 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 355.210 0.000 355.490 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 385.570 0.000 385.850 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.750 0.000 401.030 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.930 0.000 416.210 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.110 0.000 431.390 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.290 0.000 446.570 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.470 0.000 461.750 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.650 0.000 476.930 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.830 0.000 492.110 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.010 0.000 507.290 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.190 0.000 522.470 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.370 0.000 537.650 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.550 0.000 552.830 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.730 0.000 568.010 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.910 0.000 583.190 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.090 0.000 598.370 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 178.110 0.000 178.390 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 613.270 0.000 613.550 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.450 0.000 628.730 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 198.350 0.000 198.630 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 218.590 0.000 218.870 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 233.770 0.000 234.050 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 248.950 0.000 249.230 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 279.310 0.000 279.590 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 294.490 0.000 294.770 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 314.730 0.000 315.010 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 329.910 0.000 330.190 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 345.090 0.000 345.370 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 360.270 0.000 360.550 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 375.450 0.000 375.730 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 390.630 0.000 390.910 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 0.000 406.090 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.990 0.000 421.270 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.170 0.000 436.450 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.350 0.000 451.630 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 162.930 0.000 163.210 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.530 0.000 466.810 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.710 0.000 481.990 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.890 0.000 497.170 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.070 0.000 512.350 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.250 0.000 527.530 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.430 0.000 542.710 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.610 0.000 557.890 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.790 0.000 573.070 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.970 0.000 588.250 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.150 0.000 603.430 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 183.170 0.000 183.450 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.330 0.000 618.610 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.510 0.000 633.790 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 203.410 0.000 203.690 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 223.650 0.000 223.930 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 238.830 0.000 239.110 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 254.010 0.000 254.290 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 269.190 0.000 269.470 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 284.370 0.000 284.650 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 147.750 0.000 148.030 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 167.990 0.000 168.270 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 188.230 0.000 188.510 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 208.470 0.000 208.750 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 127.510 0.000 127.790 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2694.220 1487.925 ;
      LAYER met1 ;
        RECT 4.670 4.460 2695.070 1488.080 ;
      LAYER met2 ;
        RECT 4.690 1495.720 51.790 1496.410 ;
        RECT 52.630 1495.720 151.610 1496.410 ;
        RECT 152.450 1495.720 251.430 1496.410 ;
        RECT 252.270 1495.720 351.250 1496.410 ;
        RECT 352.090 1495.720 451.070 1496.410 ;
        RECT 451.910 1495.720 550.890 1496.410 ;
        RECT 551.730 1495.720 650.710 1496.410 ;
        RECT 651.550 1495.720 750.530 1496.410 ;
        RECT 751.370 1495.720 850.350 1496.410 ;
        RECT 851.190 1495.720 950.170 1496.410 ;
        RECT 951.010 1495.720 1049.990 1496.410 ;
        RECT 1050.830 1495.720 1149.810 1496.410 ;
        RECT 1150.650 1495.720 1249.630 1496.410 ;
        RECT 1250.470 1495.720 1349.450 1496.410 ;
        RECT 1350.290 1495.720 1449.270 1496.410 ;
        RECT 1450.110 1495.720 1549.090 1496.410 ;
        RECT 1549.930 1495.720 1648.910 1496.410 ;
        RECT 1649.750 1495.720 1748.730 1496.410 ;
        RECT 1749.570 1495.720 1848.550 1496.410 ;
        RECT 1849.390 1495.720 1948.370 1496.410 ;
        RECT 1949.210 1495.720 2048.190 1496.410 ;
        RECT 2049.030 1495.720 2148.010 1496.410 ;
        RECT 2148.850 1495.720 2247.830 1496.410 ;
        RECT 2248.670 1495.720 2347.650 1496.410 ;
        RECT 2348.490 1495.720 2447.470 1496.410 ;
        RECT 2448.310 1495.720 2547.290 1496.410 ;
        RECT 2548.130 1495.720 2647.110 1496.410 ;
        RECT 2647.950 1495.720 2695.050 1496.410 ;
        RECT 4.690 4.280 2695.050 1495.720 ;
        RECT 4.690 3.670 101.930 4.280 ;
        RECT 102.770 3.670 106.990 4.280 ;
        RECT 107.830 3.670 112.050 4.280 ;
        RECT 112.890 3.670 117.110 4.280 ;
        RECT 117.950 3.670 122.170 4.280 ;
        RECT 123.010 3.670 127.230 4.280 ;
        RECT 128.070 3.670 132.290 4.280 ;
        RECT 133.130 3.670 137.350 4.280 ;
        RECT 138.190 3.670 142.410 4.280 ;
        RECT 143.250 3.670 147.470 4.280 ;
        RECT 148.310 3.670 152.530 4.280 ;
        RECT 153.370 3.670 157.590 4.280 ;
        RECT 158.430 3.670 162.650 4.280 ;
        RECT 163.490 3.670 167.710 4.280 ;
        RECT 168.550 3.670 172.770 4.280 ;
        RECT 173.610 3.670 177.830 4.280 ;
        RECT 178.670 3.670 182.890 4.280 ;
        RECT 183.730 3.670 187.950 4.280 ;
        RECT 188.790 3.670 193.010 4.280 ;
        RECT 193.850 3.670 198.070 4.280 ;
        RECT 198.910 3.670 203.130 4.280 ;
        RECT 203.970 3.670 208.190 4.280 ;
        RECT 209.030 3.670 213.250 4.280 ;
        RECT 214.090 3.670 218.310 4.280 ;
        RECT 219.150 3.670 223.370 4.280 ;
        RECT 224.210 3.670 228.430 4.280 ;
        RECT 229.270 3.670 233.490 4.280 ;
        RECT 234.330 3.670 238.550 4.280 ;
        RECT 239.390 3.670 243.610 4.280 ;
        RECT 244.450 3.670 248.670 4.280 ;
        RECT 249.510 3.670 253.730 4.280 ;
        RECT 254.570 3.670 258.790 4.280 ;
        RECT 259.630 3.670 263.850 4.280 ;
        RECT 264.690 3.670 268.910 4.280 ;
        RECT 269.750 3.670 273.970 4.280 ;
        RECT 274.810 3.670 279.030 4.280 ;
        RECT 279.870 3.670 284.090 4.280 ;
        RECT 284.930 3.670 289.150 4.280 ;
        RECT 289.990 3.670 294.210 4.280 ;
        RECT 295.050 3.670 299.270 4.280 ;
        RECT 300.110 3.670 304.330 4.280 ;
        RECT 305.170 3.670 309.390 4.280 ;
        RECT 310.230 3.670 314.450 4.280 ;
        RECT 315.290 3.670 319.510 4.280 ;
        RECT 320.350 3.670 324.570 4.280 ;
        RECT 325.410 3.670 329.630 4.280 ;
        RECT 330.470 3.670 334.690 4.280 ;
        RECT 335.530 3.670 339.750 4.280 ;
        RECT 340.590 3.670 344.810 4.280 ;
        RECT 345.650 3.670 349.870 4.280 ;
        RECT 350.710 3.670 354.930 4.280 ;
        RECT 355.770 3.670 359.990 4.280 ;
        RECT 360.830 3.670 365.050 4.280 ;
        RECT 365.890 3.670 370.110 4.280 ;
        RECT 370.950 3.670 375.170 4.280 ;
        RECT 376.010 3.670 380.230 4.280 ;
        RECT 381.070 3.670 385.290 4.280 ;
        RECT 386.130 3.670 390.350 4.280 ;
        RECT 391.190 3.670 395.410 4.280 ;
        RECT 396.250 3.670 400.470 4.280 ;
        RECT 401.310 3.670 405.530 4.280 ;
        RECT 406.370 3.670 410.590 4.280 ;
        RECT 411.430 3.670 415.650 4.280 ;
        RECT 416.490 3.670 420.710 4.280 ;
        RECT 421.550 3.670 425.770 4.280 ;
        RECT 426.610 3.670 430.830 4.280 ;
        RECT 431.670 3.670 435.890 4.280 ;
        RECT 436.730 3.670 440.950 4.280 ;
        RECT 441.790 3.670 446.010 4.280 ;
        RECT 446.850 3.670 451.070 4.280 ;
        RECT 451.910 3.670 456.130 4.280 ;
        RECT 456.970 3.670 461.190 4.280 ;
        RECT 462.030 3.670 466.250 4.280 ;
        RECT 467.090 3.670 471.310 4.280 ;
        RECT 472.150 3.670 476.370 4.280 ;
        RECT 477.210 3.670 481.430 4.280 ;
        RECT 482.270 3.670 486.490 4.280 ;
        RECT 487.330 3.670 491.550 4.280 ;
        RECT 492.390 3.670 496.610 4.280 ;
        RECT 497.450 3.670 501.670 4.280 ;
        RECT 502.510 3.670 506.730 4.280 ;
        RECT 507.570 3.670 511.790 4.280 ;
        RECT 512.630 3.670 516.850 4.280 ;
        RECT 517.690 3.670 521.910 4.280 ;
        RECT 522.750 3.670 526.970 4.280 ;
        RECT 527.810 3.670 532.030 4.280 ;
        RECT 532.870 3.670 537.090 4.280 ;
        RECT 537.930 3.670 542.150 4.280 ;
        RECT 542.990 3.670 547.210 4.280 ;
        RECT 548.050 3.670 552.270 4.280 ;
        RECT 553.110 3.670 557.330 4.280 ;
        RECT 558.170 3.670 562.390 4.280 ;
        RECT 563.230 3.670 567.450 4.280 ;
        RECT 568.290 3.670 572.510 4.280 ;
        RECT 573.350 3.670 577.570 4.280 ;
        RECT 578.410 3.670 582.630 4.280 ;
        RECT 583.470 3.670 587.690 4.280 ;
        RECT 588.530 3.670 592.750 4.280 ;
        RECT 593.590 3.670 597.810 4.280 ;
        RECT 598.650 3.670 602.870 4.280 ;
        RECT 603.710 3.670 607.930 4.280 ;
        RECT 608.770 3.670 612.990 4.280 ;
        RECT 613.830 3.670 618.050 4.280 ;
        RECT 618.890 3.670 623.110 4.280 ;
        RECT 623.950 3.670 628.170 4.280 ;
        RECT 629.010 3.670 633.230 4.280 ;
        RECT 634.070 3.670 638.290 4.280 ;
        RECT 639.130 3.670 643.350 4.280 ;
        RECT 644.190 3.670 648.410 4.280 ;
        RECT 649.250 3.670 653.470 4.280 ;
        RECT 654.310 3.670 658.530 4.280 ;
        RECT 659.370 3.670 663.590 4.280 ;
        RECT 664.430 3.670 668.650 4.280 ;
        RECT 669.490 3.670 673.710 4.280 ;
        RECT 674.550 3.670 678.770 4.280 ;
        RECT 679.610 3.670 683.830 4.280 ;
        RECT 684.670 3.670 688.890 4.280 ;
        RECT 689.730 3.670 693.950 4.280 ;
        RECT 694.790 3.670 699.010 4.280 ;
        RECT 699.850 3.670 704.070 4.280 ;
        RECT 704.910 3.670 709.130 4.280 ;
        RECT 709.970 3.670 714.190 4.280 ;
        RECT 715.030 3.670 719.250 4.280 ;
        RECT 720.090 3.670 724.310 4.280 ;
        RECT 725.150 3.670 729.370 4.280 ;
        RECT 730.210 3.670 734.430 4.280 ;
        RECT 735.270 3.670 739.490 4.280 ;
        RECT 740.330 3.670 744.550 4.280 ;
        RECT 745.390 3.670 749.610 4.280 ;
        RECT 750.450 3.670 754.670 4.280 ;
        RECT 755.510 3.670 759.730 4.280 ;
        RECT 760.570 3.670 764.790 4.280 ;
        RECT 765.630 3.670 769.850 4.280 ;
        RECT 770.690 3.670 774.910 4.280 ;
        RECT 775.750 3.670 779.970 4.280 ;
        RECT 780.810 3.670 785.030 4.280 ;
        RECT 785.870 3.670 790.090 4.280 ;
        RECT 790.930 3.670 795.150 4.280 ;
        RECT 795.990 3.670 800.210 4.280 ;
        RECT 801.050 3.670 805.270 4.280 ;
        RECT 806.110 3.670 810.330 4.280 ;
        RECT 811.170 3.670 815.390 4.280 ;
        RECT 816.230 3.670 820.450 4.280 ;
        RECT 821.290 3.670 825.510 4.280 ;
        RECT 826.350 3.670 830.570 4.280 ;
        RECT 831.410 3.670 835.630 4.280 ;
        RECT 836.470 3.670 840.690 4.280 ;
        RECT 841.530 3.670 845.750 4.280 ;
        RECT 846.590 3.670 850.810 4.280 ;
        RECT 851.650 3.670 855.870 4.280 ;
        RECT 856.710 3.670 860.930 4.280 ;
        RECT 861.770 3.670 865.990 4.280 ;
        RECT 866.830 3.670 871.050 4.280 ;
        RECT 871.890 3.670 876.110 4.280 ;
        RECT 876.950 3.670 881.170 4.280 ;
        RECT 882.010 3.670 886.230 4.280 ;
        RECT 887.070 3.670 891.290 4.280 ;
        RECT 892.130 3.670 896.350 4.280 ;
        RECT 897.190 3.670 901.410 4.280 ;
        RECT 902.250 3.670 906.470 4.280 ;
        RECT 907.310 3.670 911.530 4.280 ;
        RECT 912.370 3.670 916.590 4.280 ;
        RECT 917.430 3.670 921.650 4.280 ;
        RECT 922.490 3.670 926.710 4.280 ;
        RECT 927.550 3.670 931.770 4.280 ;
        RECT 932.610 3.670 936.830 4.280 ;
        RECT 937.670 3.670 941.890 4.280 ;
        RECT 942.730 3.670 946.950 4.280 ;
        RECT 947.790 3.670 952.010 4.280 ;
        RECT 952.850 3.670 957.070 4.280 ;
        RECT 957.910 3.670 962.130 4.280 ;
        RECT 962.970 3.670 967.190 4.280 ;
        RECT 968.030 3.670 972.250 4.280 ;
        RECT 973.090 3.670 977.310 4.280 ;
        RECT 978.150 3.670 982.370 4.280 ;
        RECT 983.210 3.670 987.430 4.280 ;
        RECT 988.270 3.670 992.490 4.280 ;
        RECT 993.330 3.670 997.550 4.280 ;
        RECT 998.390 3.670 1002.610 4.280 ;
        RECT 1003.450 3.670 1007.670 4.280 ;
        RECT 1008.510 3.670 1012.730 4.280 ;
        RECT 1013.570 3.670 1017.790 4.280 ;
        RECT 1018.630 3.670 1022.850 4.280 ;
        RECT 1023.690 3.670 1027.910 4.280 ;
        RECT 1028.750 3.670 1032.970 4.280 ;
        RECT 1033.810 3.670 1038.030 4.280 ;
        RECT 1038.870 3.670 1043.090 4.280 ;
        RECT 1043.930 3.670 1048.150 4.280 ;
        RECT 1048.990 3.670 1053.210 4.280 ;
        RECT 1054.050 3.670 1058.270 4.280 ;
        RECT 1059.110 3.670 1063.330 4.280 ;
        RECT 1064.170 3.670 1068.390 4.280 ;
        RECT 1069.230 3.670 1073.450 4.280 ;
        RECT 1074.290 3.670 1078.510 4.280 ;
        RECT 1079.350 3.670 1083.570 4.280 ;
        RECT 1084.410 3.670 1088.630 4.280 ;
        RECT 1089.470 3.670 1093.690 4.280 ;
        RECT 1094.530 3.670 1098.750 4.280 ;
        RECT 1099.590 3.670 1103.810 4.280 ;
        RECT 1104.650 3.670 1108.870 4.280 ;
        RECT 1109.710 3.670 1113.930 4.280 ;
        RECT 1114.770 3.670 1118.990 4.280 ;
        RECT 1119.830 3.670 1124.050 4.280 ;
        RECT 1124.890 3.670 1129.110 4.280 ;
        RECT 1129.950 3.670 1134.170 4.280 ;
        RECT 1135.010 3.670 1139.230 4.280 ;
        RECT 1140.070 3.670 1144.290 4.280 ;
        RECT 1145.130 3.670 1149.350 4.280 ;
        RECT 1150.190 3.670 1154.410 4.280 ;
        RECT 1155.250 3.670 1159.470 4.280 ;
        RECT 1160.310 3.670 1164.530 4.280 ;
        RECT 1165.370 3.670 1169.590 4.280 ;
        RECT 1170.430 3.670 1174.650 4.280 ;
        RECT 1175.490 3.670 1179.710 4.280 ;
        RECT 1180.550 3.670 1184.770 4.280 ;
        RECT 1185.610 3.670 1189.830 4.280 ;
        RECT 1190.670 3.670 1194.890 4.280 ;
        RECT 1195.730 3.670 1199.950 4.280 ;
        RECT 1200.790 3.670 1205.010 4.280 ;
        RECT 1205.850 3.670 1210.070 4.280 ;
        RECT 1210.910 3.670 1215.130 4.280 ;
        RECT 1215.970 3.670 1220.190 4.280 ;
        RECT 1221.030 3.670 1225.250 4.280 ;
        RECT 1226.090 3.670 1230.310 4.280 ;
        RECT 1231.150 3.670 1235.370 4.280 ;
        RECT 1236.210 3.670 1240.430 4.280 ;
        RECT 1241.270 3.670 1245.490 4.280 ;
        RECT 1246.330 3.670 1250.550 4.280 ;
        RECT 1251.390 3.670 1255.610 4.280 ;
        RECT 1256.450 3.670 1260.670 4.280 ;
        RECT 1261.510 3.670 1265.730 4.280 ;
        RECT 1266.570 3.670 1270.790 4.280 ;
        RECT 1271.630 3.670 1275.850 4.280 ;
        RECT 1276.690 3.670 1280.910 4.280 ;
        RECT 1281.750 3.670 1285.970 4.280 ;
        RECT 1286.810 3.670 1291.030 4.280 ;
        RECT 1291.870 3.670 1296.090 4.280 ;
        RECT 1296.930 3.670 1301.150 4.280 ;
        RECT 1301.990 3.670 1306.210 4.280 ;
        RECT 1307.050 3.670 1311.270 4.280 ;
        RECT 1312.110 3.670 1316.330 4.280 ;
        RECT 1317.170 3.670 1321.390 4.280 ;
        RECT 1322.230 3.670 1326.450 4.280 ;
        RECT 1327.290 3.670 1331.510 4.280 ;
        RECT 1332.350 3.670 1336.570 4.280 ;
        RECT 1337.410 3.670 1341.630 4.280 ;
        RECT 1342.470 3.670 1346.690 4.280 ;
        RECT 1347.530 3.670 1351.750 4.280 ;
        RECT 1352.590 3.670 1356.810 4.280 ;
        RECT 1357.650 3.670 1361.870 4.280 ;
        RECT 1362.710 3.670 1366.930 4.280 ;
        RECT 1367.770 3.670 1371.990 4.280 ;
        RECT 1372.830 3.670 1377.050 4.280 ;
        RECT 1377.890 3.670 1382.110 4.280 ;
        RECT 1382.950 3.670 1387.170 4.280 ;
        RECT 1388.010 3.670 1392.230 4.280 ;
        RECT 1393.070 3.670 1397.290 4.280 ;
        RECT 1398.130 3.670 1402.350 4.280 ;
        RECT 1403.190 3.670 1407.410 4.280 ;
        RECT 1408.250 3.670 1412.470 4.280 ;
        RECT 1413.310 3.670 1417.530 4.280 ;
        RECT 1418.370 3.670 1422.590 4.280 ;
        RECT 1423.430 3.670 1427.650 4.280 ;
        RECT 1428.490 3.670 1432.710 4.280 ;
        RECT 1433.550 3.670 1437.770 4.280 ;
        RECT 1438.610 3.670 1442.830 4.280 ;
        RECT 1443.670 3.670 1447.890 4.280 ;
        RECT 1448.730 3.670 1452.950 4.280 ;
        RECT 1453.790 3.670 1458.010 4.280 ;
        RECT 1458.850 3.670 1463.070 4.280 ;
        RECT 1463.910 3.670 1468.130 4.280 ;
        RECT 1468.970 3.670 1473.190 4.280 ;
        RECT 1474.030 3.670 1478.250 4.280 ;
        RECT 1479.090 3.670 1483.310 4.280 ;
        RECT 1484.150 3.670 1488.370 4.280 ;
        RECT 1489.210 3.670 1493.430 4.280 ;
        RECT 1494.270 3.670 1498.490 4.280 ;
        RECT 1499.330 3.670 1503.550 4.280 ;
        RECT 1504.390 3.670 1508.610 4.280 ;
        RECT 1509.450 3.670 1513.670 4.280 ;
        RECT 1514.510 3.670 1518.730 4.280 ;
        RECT 1519.570 3.670 1523.790 4.280 ;
        RECT 1524.630 3.670 1528.850 4.280 ;
        RECT 1529.690 3.670 1533.910 4.280 ;
        RECT 1534.750 3.670 1538.970 4.280 ;
        RECT 1539.810 3.670 1544.030 4.280 ;
        RECT 1544.870 3.670 1549.090 4.280 ;
        RECT 1549.930 3.670 1554.150 4.280 ;
        RECT 1554.990 3.670 1559.210 4.280 ;
        RECT 1560.050 3.670 1564.270 4.280 ;
        RECT 1565.110 3.670 1569.330 4.280 ;
        RECT 1570.170 3.670 1574.390 4.280 ;
        RECT 1575.230 3.670 1579.450 4.280 ;
        RECT 1580.290 3.670 1584.510 4.280 ;
        RECT 1585.350 3.670 1589.570 4.280 ;
        RECT 1590.410 3.670 1594.630 4.280 ;
        RECT 1595.470 3.670 1599.690 4.280 ;
        RECT 1600.530 3.670 1604.750 4.280 ;
        RECT 1605.590 3.670 1609.810 4.280 ;
        RECT 1610.650 3.670 1614.870 4.280 ;
        RECT 1615.710 3.670 1619.930 4.280 ;
        RECT 1620.770 3.670 1624.990 4.280 ;
        RECT 1625.830 3.670 1630.050 4.280 ;
        RECT 1630.890 3.670 1635.110 4.280 ;
        RECT 1635.950 3.670 1640.170 4.280 ;
        RECT 1641.010 3.670 1645.230 4.280 ;
        RECT 1646.070 3.670 1650.290 4.280 ;
        RECT 1651.130 3.670 1655.350 4.280 ;
        RECT 1656.190 3.670 1660.410 4.280 ;
        RECT 1661.250 3.670 1665.470 4.280 ;
        RECT 1666.310 3.670 1670.530 4.280 ;
        RECT 1671.370 3.670 1675.590 4.280 ;
        RECT 1676.430 3.670 1680.650 4.280 ;
        RECT 1681.490 3.670 1685.710 4.280 ;
        RECT 1686.550 3.670 1690.770 4.280 ;
        RECT 1691.610 3.670 1695.830 4.280 ;
        RECT 1696.670 3.670 1700.890 4.280 ;
        RECT 1701.730 3.670 1705.950 4.280 ;
        RECT 1706.790 3.670 1711.010 4.280 ;
        RECT 1711.850 3.670 1716.070 4.280 ;
        RECT 1716.910 3.670 1721.130 4.280 ;
        RECT 1721.970 3.670 1726.190 4.280 ;
        RECT 1727.030 3.670 1731.250 4.280 ;
        RECT 1732.090 3.670 1736.310 4.280 ;
        RECT 1737.150 3.670 1741.370 4.280 ;
        RECT 1742.210 3.670 1746.430 4.280 ;
        RECT 1747.270 3.670 1751.490 4.280 ;
        RECT 1752.330 3.670 1756.550 4.280 ;
        RECT 1757.390 3.670 1761.610 4.280 ;
        RECT 1762.450 3.670 1766.670 4.280 ;
        RECT 1767.510 3.670 1771.730 4.280 ;
        RECT 1772.570 3.670 1776.790 4.280 ;
        RECT 1777.630 3.670 1781.850 4.280 ;
        RECT 1782.690 3.670 1786.910 4.280 ;
        RECT 1787.750 3.670 1791.970 4.280 ;
        RECT 1792.810 3.670 1797.030 4.280 ;
        RECT 1797.870 3.670 1802.090 4.280 ;
        RECT 1802.930 3.670 1807.150 4.280 ;
        RECT 1807.990 3.670 1812.210 4.280 ;
        RECT 1813.050 3.670 1817.270 4.280 ;
        RECT 1818.110 3.670 1822.330 4.280 ;
        RECT 1823.170 3.670 1827.390 4.280 ;
        RECT 1828.230 3.670 1832.450 4.280 ;
        RECT 1833.290 3.670 1837.510 4.280 ;
        RECT 1838.350 3.670 1842.570 4.280 ;
        RECT 1843.410 3.670 1847.630 4.280 ;
        RECT 1848.470 3.670 1852.690 4.280 ;
        RECT 1853.530 3.670 1857.750 4.280 ;
        RECT 1858.590 3.670 1862.810 4.280 ;
        RECT 1863.650 3.670 1867.870 4.280 ;
        RECT 1868.710 3.670 1872.930 4.280 ;
        RECT 1873.770 3.670 1877.990 4.280 ;
        RECT 1878.830 3.670 1883.050 4.280 ;
        RECT 1883.890 3.670 1888.110 4.280 ;
        RECT 1888.950 3.670 1893.170 4.280 ;
        RECT 1894.010 3.670 1898.230 4.280 ;
        RECT 1899.070 3.670 1903.290 4.280 ;
        RECT 1904.130 3.670 1908.350 4.280 ;
        RECT 1909.190 3.670 1913.410 4.280 ;
        RECT 1914.250 3.670 1918.470 4.280 ;
        RECT 1919.310 3.670 1923.530 4.280 ;
        RECT 1924.370 3.670 1928.590 4.280 ;
        RECT 1929.430 3.670 1933.650 4.280 ;
        RECT 1934.490 3.670 1938.710 4.280 ;
        RECT 1939.550 3.670 1943.770 4.280 ;
        RECT 1944.610 3.670 1948.830 4.280 ;
        RECT 1949.670 3.670 1953.890 4.280 ;
        RECT 1954.730 3.670 1958.950 4.280 ;
        RECT 1959.790 3.670 1964.010 4.280 ;
        RECT 1964.850 3.670 1969.070 4.280 ;
        RECT 1969.910 3.670 1974.130 4.280 ;
        RECT 1974.970 3.670 1979.190 4.280 ;
        RECT 1980.030 3.670 1984.250 4.280 ;
        RECT 1985.090 3.670 1989.310 4.280 ;
        RECT 1990.150 3.670 1994.370 4.280 ;
        RECT 1995.210 3.670 1999.430 4.280 ;
        RECT 2000.270 3.670 2004.490 4.280 ;
        RECT 2005.330 3.670 2009.550 4.280 ;
        RECT 2010.390 3.670 2014.610 4.280 ;
        RECT 2015.450 3.670 2019.670 4.280 ;
        RECT 2020.510 3.670 2024.730 4.280 ;
        RECT 2025.570 3.670 2029.790 4.280 ;
        RECT 2030.630 3.670 2034.850 4.280 ;
        RECT 2035.690 3.670 2039.910 4.280 ;
        RECT 2040.750 3.670 2044.970 4.280 ;
        RECT 2045.810 3.670 2050.030 4.280 ;
        RECT 2050.870 3.670 2055.090 4.280 ;
        RECT 2055.930 3.670 2060.150 4.280 ;
        RECT 2060.990 3.670 2065.210 4.280 ;
        RECT 2066.050 3.670 2070.270 4.280 ;
        RECT 2071.110 3.670 2075.330 4.280 ;
        RECT 2076.170 3.670 2080.390 4.280 ;
        RECT 2081.230 3.670 2085.450 4.280 ;
        RECT 2086.290 3.670 2090.510 4.280 ;
        RECT 2091.350 3.670 2095.570 4.280 ;
        RECT 2096.410 3.670 2100.630 4.280 ;
        RECT 2101.470 3.670 2105.690 4.280 ;
        RECT 2106.530 3.670 2110.750 4.280 ;
        RECT 2111.590 3.670 2115.810 4.280 ;
        RECT 2116.650 3.670 2120.870 4.280 ;
        RECT 2121.710 3.670 2125.930 4.280 ;
        RECT 2126.770 3.670 2130.990 4.280 ;
        RECT 2131.830 3.670 2136.050 4.280 ;
        RECT 2136.890 3.670 2141.110 4.280 ;
        RECT 2141.950 3.670 2146.170 4.280 ;
        RECT 2147.010 3.670 2151.230 4.280 ;
        RECT 2152.070 3.670 2156.290 4.280 ;
        RECT 2157.130 3.670 2161.350 4.280 ;
        RECT 2162.190 3.670 2166.410 4.280 ;
        RECT 2167.250 3.670 2171.470 4.280 ;
        RECT 2172.310 3.670 2176.530 4.280 ;
        RECT 2177.370 3.670 2181.590 4.280 ;
        RECT 2182.430 3.670 2186.650 4.280 ;
        RECT 2187.490 3.670 2191.710 4.280 ;
        RECT 2192.550 3.670 2196.770 4.280 ;
        RECT 2197.610 3.670 2201.830 4.280 ;
        RECT 2202.670 3.670 2206.890 4.280 ;
        RECT 2207.730 3.670 2211.950 4.280 ;
        RECT 2212.790 3.670 2217.010 4.280 ;
        RECT 2217.850 3.670 2222.070 4.280 ;
        RECT 2222.910 3.670 2227.130 4.280 ;
        RECT 2227.970 3.670 2232.190 4.280 ;
        RECT 2233.030 3.670 2237.250 4.280 ;
        RECT 2238.090 3.670 2242.310 4.280 ;
        RECT 2243.150 3.670 2247.370 4.280 ;
        RECT 2248.210 3.670 2252.430 4.280 ;
        RECT 2253.270 3.670 2257.490 4.280 ;
        RECT 2258.330 3.670 2262.550 4.280 ;
        RECT 2263.390 3.670 2267.610 4.280 ;
        RECT 2268.450 3.670 2272.670 4.280 ;
        RECT 2273.510 3.670 2277.730 4.280 ;
        RECT 2278.570 3.670 2282.790 4.280 ;
        RECT 2283.630 3.670 2287.850 4.280 ;
        RECT 2288.690 3.670 2292.910 4.280 ;
        RECT 2293.750 3.670 2297.970 4.280 ;
        RECT 2298.810 3.670 2303.030 4.280 ;
        RECT 2303.870 3.670 2308.090 4.280 ;
        RECT 2308.930 3.670 2313.150 4.280 ;
        RECT 2313.990 3.670 2318.210 4.280 ;
        RECT 2319.050 3.670 2323.270 4.280 ;
        RECT 2324.110 3.670 2328.330 4.280 ;
        RECT 2329.170 3.670 2333.390 4.280 ;
        RECT 2334.230 3.670 2338.450 4.280 ;
        RECT 2339.290 3.670 2343.510 4.280 ;
        RECT 2344.350 3.670 2348.570 4.280 ;
        RECT 2349.410 3.670 2353.630 4.280 ;
        RECT 2354.470 3.670 2358.690 4.280 ;
        RECT 2359.530 3.670 2363.750 4.280 ;
        RECT 2364.590 3.670 2368.810 4.280 ;
        RECT 2369.650 3.670 2373.870 4.280 ;
        RECT 2374.710 3.670 2378.930 4.280 ;
        RECT 2379.770 3.670 2383.990 4.280 ;
        RECT 2384.830 3.670 2389.050 4.280 ;
        RECT 2389.890 3.670 2394.110 4.280 ;
        RECT 2394.950 3.670 2399.170 4.280 ;
        RECT 2400.010 3.670 2404.230 4.280 ;
        RECT 2405.070 3.670 2409.290 4.280 ;
        RECT 2410.130 3.670 2414.350 4.280 ;
        RECT 2415.190 3.670 2419.410 4.280 ;
        RECT 2420.250 3.670 2424.470 4.280 ;
        RECT 2425.310 3.670 2429.530 4.280 ;
        RECT 2430.370 3.670 2434.590 4.280 ;
        RECT 2435.430 3.670 2439.650 4.280 ;
        RECT 2440.490 3.670 2444.710 4.280 ;
        RECT 2445.550 3.670 2449.770 4.280 ;
        RECT 2450.610 3.670 2454.830 4.280 ;
        RECT 2455.670 3.670 2459.890 4.280 ;
        RECT 2460.730 3.670 2464.950 4.280 ;
        RECT 2465.790 3.670 2470.010 4.280 ;
        RECT 2470.850 3.670 2475.070 4.280 ;
        RECT 2475.910 3.670 2480.130 4.280 ;
        RECT 2480.970 3.670 2485.190 4.280 ;
        RECT 2486.030 3.670 2490.250 4.280 ;
        RECT 2491.090 3.670 2495.310 4.280 ;
        RECT 2496.150 3.670 2500.370 4.280 ;
        RECT 2501.210 3.670 2505.430 4.280 ;
        RECT 2506.270 3.670 2510.490 4.280 ;
        RECT 2511.330 3.670 2515.550 4.280 ;
        RECT 2516.390 3.670 2520.610 4.280 ;
        RECT 2521.450 3.670 2525.670 4.280 ;
        RECT 2526.510 3.670 2530.730 4.280 ;
        RECT 2531.570 3.670 2535.790 4.280 ;
        RECT 2536.630 3.670 2540.850 4.280 ;
        RECT 2541.690 3.670 2545.910 4.280 ;
        RECT 2546.750 3.670 2550.970 4.280 ;
        RECT 2551.810 3.670 2556.030 4.280 ;
        RECT 2556.870 3.670 2561.090 4.280 ;
        RECT 2561.930 3.670 2566.150 4.280 ;
        RECT 2566.990 3.670 2571.210 4.280 ;
        RECT 2572.050 3.670 2576.270 4.280 ;
        RECT 2577.110 3.670 2581.330 4.280 ;
        RECT 2582.170 3.670 2586.390 4.280 ;
        RECT 2587.230 3.670 2591.450 4.280 ;
        RECT 2592.290 3.670 2596.510 4.280 ;
        RECT 2597.350 3.670 2695.050 4.280 ;
      LAYER met3 ;
        RECT 3.990 1475.280 2696.000 1488.005 ;
        RECT 4.400 1473.880 2696.000 1475.280 ;
        RECT 3.990 1468.480 2696.000 1473.880 ;
        RECT 3.990 1467.080 2695.600 1468.480 ;
        RECT 3.990 1439.920 2696.000 1467.080 ;
        RECT 4.400 1438.520 2696.000 1439.920 ;
        RECT 3.990 1435.840 2696.000 1438.520 ;
        RECT 3.990 1434.440 2695.600 1435.840 ;
        RECT 3.990 1404.560 2696.000 1434.440 ;
        RECT 4.400 1403.200 2696.000 1404.560 ;
        RECT 4.400 1403.160 2695.600 1403.200 ;
        RECT 3.990 1401.800 2695.600 1403.160 ;
        RECT 3.990 1370.560 2696.000 1401.800 ;
        RECT 3.990 1369.200 2695.600 1370.560 ;
        RECT 4.400 1369.160 2695.600 1369.200 ;
        RECT 4.400 1367.800 2696.000 1369.160 ;
        RECT 3.990 1337.920 2696.000 1367.800 ;
        RECT 3.990 1336.520 2695.600 1337.920 ;
        RECT 3.990 1333.840 2696.000 1336.520 ;
        RECT 4.400 1332.440 2696.000 1333.840 ;
        RECT 3.990 1305.280 2696.000 1332.440 ;
        RECT 3.990 1303.880 2695.600 1305.280 ;
        RECT 3.990 1298.480 2696.000 1303.880 ;
        RECT 4.400 1297.080 2696.000 1298.480 ;
        RECT 3.990 1272.640 2696.000 1297.080 ;
        RECT 3.990 1271.240 2695.600 1272.640 ;
        RECT 3.990 1263.120 2696.000 1271.240 ;
        RECT 4.400 1261.720 2696.000 1263.120 ;
        RECT 3.990 1240.000 2696.000 1261.720 ;
        RECT 3.990 1238.600 2695.600 1240.000 ;
        RECT 3.990 1227.760 2696.000 1238.600 ;
        RECT 4.400 1226.360 2696.000 1227.760 ;
        RECT 3.990 1207.360 2696.000 1226.360 ;
        RECT 3.990 1205.960 2695.600 1207.360 ;
        RECT 3.990 1192.400 2696.000 1205.960 ;
        RECT 4.400 1191.000 2696.000 1192.400 ;
        RECT 3.990 1174.720 2696.000 1191.000 ;
        RECT 3.990 1173.320 2695.600 1174.720 ;
        RECT 3.990 1157.040 2696.000 1173.320 ;
        RECT 4.400 1155.640 2696.000 1157.040 ;
        RECT 3.990 1142.080 2696.000 1155.640 ;
        RECT 3.990 1140.680 2695.600 1142.080 ;
        RECT 3.990 1121.680 2696.000 1140.680 ;
        RECT 4.400 1120.280 2696.000 1121.680 ;
        RECT 3.990 1109.440 2696.000 1120.280 ;
        RECT 3.990 1108.040 2695.600 1109.440 ;
        RECT 3.990 1086.320 2696.000 1108.040 ;
        RECT 4.400 1084.920 2696.000 1086.320 ;
        RECT 3.990 1076.800 2696.000 1084.920 ;
        RECT 3.990 1075.400 2695.600 1076.800 ;
        RECT 3.990 1050.960 2696.000 1075.400 ;
        RECT 4.400 1049.560 2696.000 1050.960 ;
        RECT 3.990 1044.160 2696.000 1049.560 ;
        RECT 3.990 1042.760 2695.600 1044.160 ;
        RECT 3.990 1015.600 2696.000 1042.760 ;
        RECT 4.400 1014.200 2696.000 1015.600 ;
        RECT 3.990 1011.520 2696.000 1014.200 ;
        RECT 3.990 1010.120 2695.600 1011.520 ;
        RECT 3.990 980.240 2696.000 1010.120 ;
        RECT 4.400 978.880 2696.000 980.240 ;
        RECT 4.400 978.840 2695.600 978.880 ;
        RECT 3.990 977.480 2695.600 978.840 ;
        RECT 3.990 946.240 2696.000 977.480 ;
        RECT 3.990 944.880 2695.600 946.240 ;
        RECT 4.400 944.840 2695.600 944.880 ;
        RECT 4.400 943.480 2696.000 944.840 ;
        RECT 3.990 913.600 2696.000 943.480 ;
        RECT 3.990 912.200 2695.600 913.600 ;
        RECT 3.990 909.520 2696.000 912.200 ;
        RECT 4.400 908.120 2696.000 909.520 ;
        RECT 3.990 880.960 2696.000 908.120 ;
        RECT 3.990 879.560 2695.600 880.960 ;
        RECT 3.990 874.160 2696.000 879.560 ;
        RECT 4.400 872.760 2696.000 874.160 ;
        RECT 3.990 848.320 2696.000 872.760 ;
        RECT 3.990 846.920 2695.600 848.320 ;
        RECT 3.990 838.800 2696.000 846.920 ;
        RECT 4.400 837.400 2696.000 838.800 ;
        RECT 3.990 815.680 2696.000 837.400 ;
        RECT 3.990 814.280 2695.600 815.680 ;
        RECT 3.990 803.440 2696.000 814.280 ;
        RECT 4.400 802.040 2696.000 803.440 ;
        RECT 3.990 783.040 2696.000 802.040 ;
        RECT 3.990 781.640 2695.600 783.040 ;
        RECT 3.990 768.080 2696.000 781.640 ;
        RECT 4.400 766.680 2696.000 768.080 ;
        RECT 3.990 750.400 2696.000 766.680 ;
        RECT 3.990 749.000 2695.600 750.400 ;
        RECT 3.990 732.720 2696.000 749.000 ;
        RECT 4.400 731.320 2696.000 732.720 ;
        RECT 3.990 717.760 2696.000 731.320 ;
        RECT 3.990 716.360 2695.600 717.760 ;
        RECT 3.990 697.360 2696.000 716.360 ;
        RECT 4.400 695.960 2696.000 697.360 ;
        RECT 3.990 685.120 2696.000 695.960 ;
        RECT 3.990 683.720 2695.600 685.120 ;
        RECT 3.990 662.000 2696.000 683.720 ;
        RECT 4.400 660.600 2696.000 662.000 ;
        RECT 3.990 652.480 2696.000 660.600 ;
        RECT 3.990 651.080 2695.600 652.480 ;
        RECT 3.990 626.640 2696.000 651.080 ;
        RECT 4.400 625.240 2696.000 626.640 ;
        RECT 3.990 619.840 2696.000 625.240 ;
        RECT 3.990 618.440 2695.600 619.840 ;
        RECT 3.990 591.280 2696.000 618.440 ;
        RECT 4.400 589.880 2696.000 591.280 ;
        RECT 3.990 587.200 2696.000 589.880 ;
        RECT 3.990 585.800 2695.600 587.200 ;
        RECT 3.990 555.920 2696.000 585.800 ;
        RECT 4.400 554.560 2696.000 555.920 ;
        RECT 4.400 554.520 2695.600 554.560 ;
        RECT 3.990 553.160 2695.600 554.520 ;
        RECT 3.990 521.920 2696.000 553.160 ;
        RECT 3.990 520.560 2695.600 521.920 ;
        RECT 4.400 520.520 2695.600 520.560 ;
        RECT 4.400 519.160 2696.000 520.520 ;
        RECT 3.990 489.280 2696.000 519.160 ;
        RECT 3.990 487.880 2695.600 489.280 ;
        RECT 3.990 485.200 2696.000 487.880 ;
        RECT 4.400 483.800 2696.000 485.200 ;
        RECT 3.990 456.640 2696.000 483.800 ;
        RECT 3.990 455.240 2695.600 456.640 ;
        RECT 3.990 449.840 2696.000 455.240 ;
        RECT 4.400 448.440 2696.000 449.840 ;
        RECT 3.990 424.000 2696.000 448.440 ;
        RECT 3.990 422.600 2695.600 424.000 ;
        RECT 3.990 414.480 2696.000 422.600 ;
        RECT 4.400 413.080 2696.000 414.480 ;
        RECT 3.990 391.360 2696.000 413.080 ;
        RECT 3.990 389.960 2695.600 391.360 ;
        RECT 3.990 379.120 2696.000 389.960 ;
        RECT 4.400 377.720 2696.000 379.120 ;
        RECT 3.990 358.720 2696.000 377.720 ;
        RECT 3.990 357.320 2695.600 358.720 ;
        RECT 3.990 343.760 2696.000 357.320 ;
        RECT 4.400 342.360 2696.000 343.760 ;
        RECT 3.990 326.080 2696.000 342.360 ;
        RECT 3.990 324.680 2695.600 326.080 ;
        RECT 3.990 308.400 2696.000 324.680 ;
        RECT 4.400 307.000 2696.000 308.400 ;
        RECT 3.990 293.440 2696.000 307.000 ;
        RECT 3.990 292.040 2695.600 293.440 ;
        RECT 3.990 273.040 2696.000 292.040 ;
        RECT 4.400 271.640 2696.000 273.040 ;
        RECT 3.990 260.800 2696.000 271.640 ;
        RECT 3.990 259.400 2695.600 260.800 ;
        RECT 3.990 237.680 2696.000 259.400 ;
        RECT 4.400 236.280 2696.000 237.680 ;
        RECT 3.990 228.160 2696.000 236.280 ;
        RECT 3.990 226.760 2695.600 228.160 ;
        RECT 3.990 202.320 2696.000 226.760 ;
        RECT 4.400 200.920 2696.000 202.320 ;
        RECT 3.990 195.520 2696.000 200.920 ;
        RECT 3.990 194.120 2695.600 195.520 ;
        RECT 3.990 166.960 2696.000 194.120 ;
        RECT 4.400 165.560 2696.000 166.960 ;
        RECT 3.990 162.880 2696.000 165.560 ;
        RECT 3.990 161.480 2695.600 162.880 ;
        RECT 3.990 131.600 2696.000 161.480 ;
        RECT 4.400 130.240 2696.000 131.600 ;
        RECT 4.400 130.200 2695.600 130.240 ;
        RECT 3.990 128.840 2695.600 130.200 ;
        RECT 3.990 97.600 2696.000 128.840 ;
        RECT 3.990 96.240 2695.600 97.600 ;
        RECT 4.400 96.200 2695.600 96.240 ;
        RECT 4.400 94.840 2696.000 96.200 ;
        RECT 3.990 64.960 2696.000 94.840 ;
        RECT 3.990 63.560 2695.600 64.960 ;
        RECT 3.990 60.880 2696.000 63.560 ;
        RECT 4.400 59.480 2696.000 60.880 ;
        RECT 3.990 32.320 2696.000 59.480 ;
        RECT 3.990 30.920 2695.600 32.320 ;
        RECT 3.990 25.520 2696.000 30.920 ;
        RECT 4.400 24.120 2696.000 25.520 ;
        RECT 3.990 6.295 2696.000 24.120 ;
      LAYER met4 ;
        RECT 1544.975 194.655 1556.640 396.945 ;
        RECT 1559.040 194.655 1633.440 396.945 ;
        RECT 1635.840 194.655 1710.240 396.945 ;
        RECT 1712.640 194.655 1787.040 396.945 ;
        RECT 1789.440 194.655 1863.840 396.945 ;
        RECT 1866.240 194.655 1940.640 396.945 ;
        RECT 1943.040 194.655 2017.440 396.945 ;
        RECT 2019.840 194.655 2076.145 396.945 ;
  END
END user_proj_example
END LIBRARY

