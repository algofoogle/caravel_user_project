magic
tech sky130A
magscale 1 2
timestamp 1727304141
<< obsli1 >>
rect 1104 2159 538844 297585
<< obsm1 >>
rect 934 892 539014 297616
<< metal2 >>
rect 10414 299200 10470 300000
rect 30378 299200 30434 300000
rect 50342 299200 50398 300000
rect 70306 299200 70362 300000
rect 90270 299200 90326 300000
rect 110234 299200 110290 300000
rect 130198 299200 130254 300000
rect 150162 299200 150218 300000
rect 170126 299200 170182 300000
rect 190090 299200 190146 300000
rect 210054 299200 210110 300000
rect 230018 299200 230074 300000
rect 249982 299200 250038 300000
rect 269946 299200 270002 300000
rect 289910 299200 289966 300000
rect 309874 299200 309930 300000
rect 329838 299200 329894 300000
rect 349802 299200 349858 300000
rect 369766 299200 369822 300000
rect 389730 299200 389786 300000
rect 409694 299200 409750 300000
rect 429658 299200 429714 300000
rect 449622 299200 449678 300000
rect 469586 299200 469642 300000
rect 489550 299200 489606 300000
rect 509514 299200 509570 300000
rect 529478 299200 529534 300000
rect 20442 0 20498 800
rect 21454 0 21510 800
rect 22466 0 22522 800
rect 23478 0 23534 800
rect 24490 0 24546 800
rect 25502 0 25558 800
rect 26514 0 26570 800
rect 27526 0 27582 800
rect 28538 0 28594 800
rect 29550 0 29606 800
rect 30562 0 30618 800
rect 31574 0 31630 800
rect 32586 0 32642 800
rect 33598 0 33654 800
rect 34610 0 34666 800
rect 35622 0 35678 800
rect 36634 0 36690 800
rect 37646 0 37702 800
rect 38658 0 38714 800
rect 39670 0 39726 800
rect 40682 0 40738 800
rect 41694 0 41750 800
rect 42706 0 42762 800
rect 43718 0 43774 800
rect 44730 0 44786 800
rect 45742 0 45798 800
rect 46754 0 46810 800
rect 47766 0 47822 800
rect 48778 0 48834 800
rect 49790 0 49846 800
rect 50802 0 50858 800
rect 51814 0 51870 800
rect 52826 0 52882 800
rect 53838 0 53894 800
rect 54850 0 54906 800
rect 55862 0 55918 800
rect 56874 0 56930 800
rect 57886 0 57942 800
rect 58898 0 58954 800
rect 59910 0 59966 800
rect 60922 0 60978 800
rect 61934 0 61990 800
rect 62946 0 63002 800
rect 63958 0 64014 800
rect 64970 0 65026 800
rect 65982 0 66038 800
rect 66994 0 67050 800
rect 68006 0 68062 800
rect 69018 0 69074 800
rect 70030 0 70086 800
rect 71042 0 71098 800
rect 72054 0 72110 800
rect 73066 0 73122 800
rect 74078 0 74134 800
rect 75090 0 75146 800
rect 76102 0 76158 800
rect 77114 0 77170 800
rect 78126 0 78182 800
rect 79138 0 79194 800
rect 80150 0 80206 800
rect 81162 0 81218 800
rect 82174 0 82230 800
rect 83186 0 83242 800
rect 84198 0 84254 800
rect 85210 0 85266 800
rect 86222 0 86278 800
rect 87234 0 87290 800
rect 88246 0 88302 800
rect 89258 0 89314 800
rect 90270 0 90326 800
rect 91282 0 91338 800
rect 92294 0 92350 800
rect 93306 0 93362 800
rect 94318 0 94374 800
rect 95330 0 95386 800
rect 96342 0 96398 800
rect 97354 0 97410 800
rect 98366 0 98422 800
rect 99378 0 99434 800
rect 100390 0 100446 800
rect 101402 0 101458 800
rect 102414 0 102470 800
rect 103426 0 103482 800
rect 104438 0 104494 800
rect 105450 0 105506 800
rect 106462 0 106518 800
rect 107474 0 107530 800
rect 108486 0 108542 800
rect 109498 0 109554 800
rect 110510 0 110566 800
rect 111522 0 111578 800
rect 112534 0 112590 800
rect 113546 0 113602 800
rect 114558 0 114614 800
rect 115570 0 115626 800
rect 116582 0 116638 800
rect 117594 0 117650 800
rect 118606 0 118662 800
rect 119618 0 119674 800
rect 120630 0 120686 800
rect 121642 0 121698 800
rect 122654 0 122710 800
rect 123666 0 123722 800
rect 124678 0 124734 800
rect 125690 0 125746 800
rect 126702 0 126758 800
rect 127714 0 127770 800
rect 128726 0 128782 800
rect 129738 0 129794 800
rect 130750 0 130806 800
rect 131762 0 131818 800
rect 132774 0 132830 800
rect 133786 0 133842 800
rect 134798 0 134854 800
rect 135810 0 135866 800
rect 136822 0 136878 800
rect 137834 0 137890 800
rect 138846 0 138902 800
rect 139858 0 139914 800
rect 140870 0 140926 800
rect 141882 0 141938 800
rect 142894 0 142950 800
rect 143906 0 143962 800
rect 144918 0 144974 800
rect 145930 0 145986 800
rect 146942 0 146998 800
rect 147954 0 148010 800
rect 148966 0 149022 800
rect 149978 0 150034 800
rect 150990 0 151046 800
rect 152002 0 152058 800
rect 153014 0 153070 800
rect 154026 0 154082 800
rect 155038 0 155094 800
rect 156050 0 156106 800
rect 157062 0 157118 800
rect 158074 0 158130 800
rect 159086 0 159142 800
rect 160098 0 160154 800
rect 161110 0 161166 800
rect 162122 0 162178 800
rect 163134 0 163190 800
rect 164146 0 164202 800
rect 165158 0 165214 800
rect 166170 0 166226 800
rect 167182 0 167238 800
rect 168194 0 168250 800
rect 169206 0 169262 800
rect 170218 0 170274 800
rect 171230 0 171286 800
rect 172242 0 172298 800
rect 173254 0 173310 800
rect 174266 0 174322 800
rect 175278 0 175334 800
rect 176290 0 176346 800
rect 177302 0 177358 800
rect 178314 0 178370 800
rect 179326 0 179382 800
rect 180338 0 180394 800
rect 181350 0 181406 800
rect 182362 0 182418 800
rect 183374 0 183430 800
rect 184386 0 184442 800
rect 185398 0 185454 800
rect 186410 0 186466 800
rect 187422 0 187478 800
rect 188434 0 188490 800
rect 189446 0 189502 800
rect 190458 0 190514 800
rect 191470 0 191526 800
rect 192482 0 192538 800
rect 193494 0 193550 800
rect 194506 0 194562 800
rect 195518 0 195574 800
rect 196530 0 196586 800
rect 197542 0 197598 800
rect 198554 0 198610 800
rect 199566 0 199622 800
rect 200578 0 200634 800
rect 201590 0 201646 800
rect 202602 0 202658 800
rect 203614 0 203670 800
rect 204626 0 204682 800
rect 205638 0 205694 800
rect 206650 0 206706 800
rect 207662 0 207718 800
rect 208674 0 208730 800
rect 209686 0 209742 800
rect 210698 0 210754 800
rect 211710 0 211766 800
rect 212722 0 212778 800
rect 213734 0 213790 800
rect 214746 0 214802 800
rect 215758 0 215814 800
rect 216770 0 216826 800
rect 217782 0 217838 800
rect 218794 0 218850 800
rect 219806 0 219862 800
rect 220818 0 220874 800
rect 221830 0 221886 800
rect 222842 0 222898 800
rect 223854 0 223910 800
rect 224866 0 224922 800
rect 225878 0 225934 800
rect 226890 0 226946 800
rect 227902 0 227958 800
rect 228914 0 228970 800
rect 229926 0 229982 800
rect 230938 0 230994 800
rect 231950 0 232006 800
rect 232962 0 233018 800
rect 233974 0 234030 800
rect 234986 0 235042 800
rect 235998 0 236054 800
rect 237010 0 237066 800
rect 238022 0 238078 800
rect 239034 0 239090 800
rect 240046 0 240102 800
rect 241058 0 241114 800
rect 242070 0 242126 800
rect 243082 0 243138 800
rect 244094 0 244150 800
rect 245106 0 245162 800
rect 246118 0 246174 800
rect 247130 0 247186 800
rect 248142 0 248198 800
rect 249154 0 249210 800
rect 250166 0 250222 800
rect 251178 0 251234 800
rect 252190 0 252246 800
rect 253202 0 253258 800
rect 254214 0 254270 800
rect 255226 0 255282 800
rect 256238 0 256294 800
rect 257250 0 257306 800
rect 258262 0 258318 800
rect 259274 0 259330 800
rect 260286 0 260342 800
rect 261298 0 261354 800
rect 262310 0 262366 800
rect 263322 0 263378 800
rect 264334 0 264390 800
rect 265346 0 265402 800
rect 266358 0 266414 800
rect 267370 0 267426 800
rect 268382 0 268438 800
rect 269394 0 269450 800
rect 270406 0 270462 800
rect 271418 0 271474 800
rect 272430 0 272486 800
rect 273442 0 273498 800
rect 274454 0 274510 800
rect 275466 0 275522 800
rect 276478 0 276534 800
rect 277490 0 277546 800
rect 278502 0 278558 800
rect 279514 0 279570 800
rect 280526 0 280582 800
rect 281538 0 281594 800
rect 282550 0 282606 800
rect 283562 0 283618 800
rect 284574 0 284630 800
rect 285586 0 285642 800
rect 286598 0 286654 800
rect 287610 0 287666 800
rect 288622 0 288678 800
rect 289634 0 289690 800
rect 290646 0 290702 800
rect 291658 0 291714 800
rect 292670 0 292726 800
rect 293682 0 293738 800
rect 294694 0 294750 800
rect 295706 0 295762 800
rect 296718 0 296774 800
rect 297730 0 297786 800
rect 298742 0 298798 800
rect 299754 0 299810 800
rect 300766 0 300822 800
rect 301778 0 301834 800
rect 302790 0 302846 800
rect 303802 0 303858 800
rect 304814 0 304870 800
rect 305826 0 305882 800
rect 306838 0 306894 800
rect 307850 0 307906 800
rect 308862 0 308918 800
rect 309874 0 309930 800
rect 310886 0 310942 800
rect 311898 0 311954 800
rect 312910 0 312966 800
rect 313922 0 313978 800
rect 314934 0 314990 800
rect 315946 0 316002 800
rect 316958 0 317014 800
rect 317970 0 318026 800
rect 318982 0 319038 800
rect 319994 0 320050 800
rect 321006 0 321062 800
rect 322018 0 322074 800
rect 323030 0 323086 800
rect 324042 0 324098 800
rect 325054 0 325110 800
rect 326066 0 326122 800
rect 327078 0 327134 800
rect 328090 0 328146 800
rect 329102 0 329158 800
rect 330114 0 330170 800
rect 331126 0 331182 800
rect 332138 0 332194 800
rect 333150 0 333206 800
rect 334162 0 334218 800
rect 335174 0 335230 800
rect 336186 0 336242 800
rect 337198 0 337254 800
rect 338210 0 338266 800
rect 339222 0 339278 800
rect 340234 0 340290 800
rect 341246 0 341302 800
rect 342258 0 342314 800
rect 343270 0 343326 800
rect 344282 0 344338 800
rect 345294 0 345350 800
rect 346306 0 346362 800
rect 347318 0 347374 800
rect 348330 0 348386 800
rect 349342 0 349398 800
rect 350354 0 350410 800
rect 351366 0 351422 800
rect 352378 0 352434 800
rect 353390 0 353446 800
rect 354402 0 354458 800
rect 355414 0 355470 800
rect 356426 0 356482 800
rect 357438 0 357494 800
rect 358450 0 358506 800
rect 359462 0 359518 800
rect 360474 0 360530 800
rect 361486 0 361542 800
rect 362498 0 362554 800
rect 363510 0 363566 800
rect 364522 0 364578 800
rect 365534 0 365590 800
rect 366546 0 366602 800
rect 367558 0 367614 800
rect 368570 0 368626 800
rect 369582 0 369638 800
rect 370594 0 370650 800
rect 371606 0 371662 800
rect 372618 0 372674 800
rect 373630 0 373686 800
rect 374642 0 374698 800
rect 375654 0 375710 800
rect 376666 0 376722 800
rect 377678 0 377734 800
rect 378690 0 378746 800
rect 379702 0 379758 800
rect 380714 0 380770 800
rect 381726 0 381782 800
rect 382738 0 382794 800
rect 383750 0 383806 800
rect 384762 0 384818 800
rect 385774 0 385830 800
rect 386786 0 386842 800
rect 387798 0 387854 800
rect 388810 0 388866 800
rect 389822 0 389878 800
rect 390834 0 390890 800
rect 391846 0 391902 800
rect 392858 0 392914 800
rect 393870 0 393926 800
rect 394882 0 394938 800
rect 395894 0 395950 800
rect 396906 0 396962 800
rect 397918 0 397974 800
rect 398930 0 398986 800
rect 399942 0 399998 800
rect 400954 0 401010 800
rect 401966 0 402022 800
rect 402978 0 403034 800
rect 403990 0 404046 800
rect 405002 0 405058 800
rect 406014 0 406070 800
rect 407026 0 407082 800
rect 408038 0 408094 800
rect 409050 0 409106 800
rect 410062 0 410118 800
rect 411074 0 411130 800
rect 412086 0 412142 800
rect 413098 0 413154 800
rect 414110 0 414166 800
rect 415122 0 415178 800
rect 416134 0 416190 800
rect 417146 0 417202 800
rect 418158 0 418214 800
rect 419170 0 419226 800
rect 420182 0 420238 800
rect 421194 0 421250 800
rect 422206 0 422262 800
rect 423218 0 423274 800
rect 424230 0 424286 800
rect 425242 0 425298 800
rect 426254 0 426310 800
rect 427266 0 427322 800
rect 428278 0 428334 800
rect 429290 0 429346 800
rect 430302 0 430358 800
rect 431314 0 431370 800
rect 432326 0 432382 800
rect 433338 0 433394 800
rect 434350 0 434406 800
rect 435362 0 435418 800
rect 436374 0 436430 800
rect 437386 0 437442 800
rect 438398 0 438454 800
rect 439410 0 439466 800
rect 440422 0 440478 800
rect 441434 0 441490 800
rect 442446 0 442502 800
rect 443458 0 443514 800
rect 444470 0 444526 800
rect 445482 0 445538 800
rect 446494 0 446550 800
rect 447506 0 447562 800
rect 448518 0 448574 800
rect 449530 0 449586 800
rect 450542 0 450598 800
rect 451554 0 451610 800
rect 452566 0 452622 800
rect 453578 0 453634 800
rect 454590 0 454646 800
rect 455602 0 455658 800
rect 456614 0 456670 800
rect 457626 0 457682 800
rect 458638 0 458694 800
rect 459650 0 459706 800
rect 460662 0 460718 800
rect 461674 0 461730 800
rect 462686 0 462742 800
rect 463698 0 463754 800
rect 464710 0 464766 800
rect 465722 0 465778 800
rect 466734 0 466790 800
rect 467746 0 467802 800
rect 468758 0 468814 800
rect 469770 0 469826 800
rect 470782 0 470838 800
rect 471794 0 471850 800
rect 472806 0 472862 800
rect 473818 0 473874 800
rect 474830 0 474886 800
rect 475842 0 475898 800
rect 476854 0 476910 800
rect 477866 0 477922 800
rect 478878 0 478934 800
rect 479890 0 479946 800
rect 480902 0 480958 800
rect 481914 0 481970 800
rect 482926 0 482982 800
rect 483938 0 483994 800
rect 484950 0 485006 800
rect 485962 0 486018 800
rect 486974 0 487030 800
rect 487986 0 488042 800
rect 488998 0 489054 800
rect 490010 0 490066 800
rect 491022 0 491078 800
rect 492034 0 492090 800
rect 493046 0 493102 800
rect 494058 0 494114 800
rect 495070 0 495126 800
rect 496082 0 496138 800
rect 497094 0 497150 800
rect 498106 0 498162 800
rect 499118 0 499174 800
rect 500130 0 500186 800
rect 501142 0 501198 800
rect 502154 0 502210 800
rect 503166 0 503222 800
rect 504178 0 504234 800
rect 505190 0 505246 800
rect 506202 0 506258 800
rect 507214 0 507270 800
rect 508226 0 508282 800
rect 509238 0 509294 800
rect 510250 0 510306 800
rect 511262 0 511318 800
rect 512274 0 512330 800
rect 513286 0 513342 800
rect 514298 0 514354 800
rect 515310 0 515366 800
rect 516322 0 516378 800
rect 517334 0 517390 800
rect 518346 0 518402 800
rect 519358 0 519414 800
<< obsm2 >>
rect 938 299144 10358 299282
rect 10526 299144 30322 299282
rect 30490 299144 50286 299282
rect 50454 299144 70250 299282
rect 70418 299144 90214 299282
rect 90382 299144 110178 299282
rect 110346 299144 130142 299282
rect 130310 299144 150106 299282
rect 150274 299144 170070 299282
rect 170238 299144 190034 299282
rect 190202 299144 209998 299282
rect 210166 299144 229962 299282
rect 230130 299144 249926 299282
rect 250094 299144 269890 299282
rect 270058 299144 289854 299282
rect 290022 299144 309818 299282
rect 309986 299144 329782 299282
rect 329950 299144 349746 299282
rect 349914 299144 369710 299282
rect 369878 299144 389674 299282
rect 389842 299144 409638 299282
rect 409806 299144 429602 299282
rect 429770 299144 449566 299282
rect 449734 299144 469530 299282
rect 469698 299144 489494 299282
rect 489662 299144 509458 299282
rect 509626 299144 529422 299282
rect 529590 299144 539010 299282
rect 938 856 539010 299144
rect 938 734 20386 856
rect 20554 734 21398 856
rect 21566 734 22410 856
rect 22578 734 23422 856
rect 23590 734 24434 856
rect 24602 734 25446 856
rect 25614 734 26458 856
rect 26626 734 27470 856
rect 27638 734 28482 856
rect 28650 734 29494 856
rect 29662 734 30506 856
rect 30674 734 31518 856
rect 31686 734 32530 856
rect 32698 734 33542 856
rect 33710 734 34554 856
rect 34722 734 35566 856
rect 35734 734 36578 856
rect 36746 734 37590 856
rect 37758 734 38602 856
rect 38770 734 39614 856
rect 39782 734 40626 856
rect 40794 734 41638 856
rect 41806 734 42650 856
rect 42818 734 43662 856
rect 43830 734 44674 856
rect 44842 734 45686 856
rect 45854 734 46698 856
rect 46866 734 47710 856
rect 47878 734 48722 856
rect 48890 734 49734 856
rect 49902 734 50746 856
rect 50914 734 51758 856
rect 51926 734 52770 856
rect 52938 734 53782 856
rect 53950 734 54794 856
rect 54962 734 55806 856
rect 55974 734 56818 856
rect 56986 734 57830 856
rect 57998 734 58842 856
rect 59010 734 59854 856
rect 60022 734 60866 856
rect 61034 734 61878 856
rect 62046 734 62890 856
rect 63058 734 63902 856
rect 64070 734 64914 856
rect 65082 734 65926 856
rect 66094 734 66938 856
rect 67106 734 67950 856
rect 68118 734 68962 856
rect 69130 734 69974 856
rect 70142 734 70986 856
rect 71154 734 71998 856
rect 72166 734 73010 856
rect 73178 734 74022 856
rect 74190 734 75034 856
rect 75202 734 76046 856
rect 76214 734 77058 856
rect 77226 734 78070 856
rect 78238 734 79082 856
rect 79250 734 80094 856
rect 80262 734 81106 856
rect 81274 734 82118 856
rect 82286 734 83130 856
rect 83298 734 84142 856
rect 84310 734 85154 856
rect 85322 734 86166 856
rect 86334 734 87178 856
rect 87346 734 88190 856
rect 88358 734 89202 856
rect 89370 734 90214 856
rect 90382 734 91226 856
rect 91394 734 92238 856
rect 92406 734 93250 856
rect 93418 734 94262 856
rect 94430 734 95274 856
rect 95442 734 96286 856
rect 96454 734 97298 856
rect 97466 734 98310 856
rect 98478 734 99322 856
rect 99490 734 100334 856
rect 100502 734 101346 856
rect 101514 734 102358 856
rect 102526 734 103370 856
rect 103538 734 104382 856
rect 104550 734 105394 856
rect 105562 734 106406 856
rect 106574 734 107418 856
rect 107586 734 108430 856
rect 108598 734 109442 856
rect 109610 734 110454 856
rect 110622 734 111466 856
rect 111634 734 112478 856
rect 112646 734 113490 856
rect 113658 734 114502 856
rect 114670 734 115514 856
rect 115682 734 116526 856
rect 116694 734 117538 856
rect 117706 734 118550 856
rect 118718 734 119562 856
rect 119730 734 120574 856
rect 120742 734 121586 856
rect 121754 734 122598 856
rect 122766 734 123610 856
rect 123778 734 124622 856
rect 124790 734 125634 856
rect 125802 734 126646 856
rect 126814 734 127658 856
rect 127826 734 128670 856
rect 128838 734 129682 856
rect 129850 734 130694 856
rect 130862 734 131706 856
rect 131874 734 132718 856
rect 132886 734 133730 856
rect 133898 734 134742 856
rect 134910 734 135754 856
rect 135922 734 136766 856
rect 136934 734 137778 856
rect 137946 734 138790 856
rect 138958 734 139802 856
rect 139970 734 140814 856
rect 140982 734 141826 856
rect 141994 734 142838 856
rect 143006 734 143850 856
rect 144018 734 144862 856
rect 145030 734 145874 856
rect 146042 734 146886 856
rect 147054 734 147898 856
rect 148066 734 148910 856
rect 149078 734 149922 856
rect 150090 734 150934 856
rect 151102 734 151946 856
rect 152114 734 152958 856
rect 153126 734 153970 856
rect 154138 734 154982 856
rect 155150 734 155994 856
rect 156162 734 157006 856
rect 157174 734 158018 856
rect 158186 734 159030 856
rect 159198 734 160042 856
rect 160210 734 161054 856
rect 161222 734 162066 856
rect 162234 734 163078 856
rect 163246 734 164090 856
rect 164258 734 165102 856
rect 165270 734 166114 856
rect 166282 734 167126 856
rect 167294 734 168138 856
rect 168306 734 169150 856
rect 169318 734 170162 856
rect 170330 734 171174 856
rect 171342 734 172186 856
rect 172354 734 173198 856
rect 173366 734 174210 856
rect 174378 734 175222 856
rect 175390 734 176234 856
rect 176402 734 177246 856
rect 177414 734 178258 856
rect 178426 734 179270 856
rect 179438 734 180282 856
rect 180450 734 181294 856
rect 181462 734 182306 856
rect 182474 734 183318 856
rect 183486 734 184330 856
rect 184498 734 185342 856
rect 185510 734 186354 856
rect 186522 734 187366 856
rect 187534 734 188378 856
rect 188546 734 189390 856
rect 189558 734 190402 856
rect 190570 734 191414 856
rect 191582 734 192426 856
rect 192594 734 193438 856
rect 193606 734 194450 856
rect 194618 734 195462 856
rect 195630 734 196474 856
rect 196642 734 197486 856
rect 197654 734 198498 856
rect 198666 734 199510 856
rect 199678 734 200522 856
rect 200690 734 201534 856
rect 201702 734 202546 856
rect 202714 734 203558 856
rect 203726 734 204570 856
rect 204738 734 205582 856
rect 205750 734 206594 856
rect 206762 734 207606 856
rect 207774 734 208618 856
rect 208786 734 209630 856
rect 209798 734 210642 856
rect 210810 734 211654 856
rect 211822 734 212666 856
rect 212834 734 213678 856
rect 213846 734 214690 856
rect 214858 734 215702 856
rect 215870 734 216714 856
rect 216882 734 217726 856
rect 217894 734 218738 856
rect 218906 734 219750 856
rect 219918 734 220762 856
rect 220930 734 221774 856
rect 221942 734 222786 856
rect 222954 734 223798 856
rect 223966 734 224810 856
rect 224978 734 225822 856
rect 225990 734 226834 856
rect 227002 734 227846 856
rect 228014 734 228858 856
rect 229026 734 229870 856
rect 230038 734 230882 856
rect 231050 734 231894 856
rect 232062 734 232906 856
rect 233074 734 233918 856
rect 234086 734 234930 856
rect 235098 734 235942 856
rect 236110 734 236954 856
rect 237122 734 237966 856
rect 238134 734 238978 856
rect 239146 734 239990 856
rect 240158 734 241002 856
rect 241170 734 242014 856
rect 242182 734 243026 856
rect 243194 734 244038 856
rect 244206 734 245050 856
rect 245218 734 246062 856
rect 246230 734 247074 856
rect 247242 734 248086 856
rect 248254 734 249098 856
rect 249266 734 250110 856
rect 250278 734 251122 856
rect 251290 734 252134 856
rect 252302 734 253146 856
rect 253314 734 254158 856
rect 254326 734 255170 856
rect 255338 734 256182 856
rect 256350 734 257194 856
rect 257362 734 258206 856
rect 258374 734 259218 856
rect 259386 734 260230 856
rect 260398 734 261242 856
rect 261410 734 262254 856
rect 262422 734 263266 856
rect 263434 734 264278 856
rect 264446 734 265290 856
rect 265458 734 266302 856
rect 266470 734 267314 856
rect 267482 734 268326 856
rect 268494 734 269338 856
rect 269506 734 270350 856
rect 270518 734 271362 856
rect 271530 734 272374 856
rect 272542 734 273386 856
rect 273554 734 274398 856
rect 274566 734 275410 856
rect 275578 734 276422 856
rect 276590 734 277434 856
rect 277602 734 278446 856
rect 278614 734 279458 856
rect 279626 734 280470 856
rect 280638 734 281482 856
rect 281650 734 282494 856
rect 282662 734 283506 856
rect 283674 734 284518 856
rect 284686 734 285530 856
rect 285698 734 286542 856
rect 286710 734 287554 856
rect 287722 734 288566 856
rect 288734 734 289578 856
rect 289746 734 290590 856
rect 290758 734 291602 856
rect 291770 734 292614 856
rect 292782 734 293626 856
rect 293794 734 294638 856
rect 294806 734 295650 856
rect 295818 734 296662 856
rect 296830 734 297674 856
rect 297842 734 298686 856
rect 298854 734 299698 856
rect 299866 734 300710 856
rect 300878 734 301722 856
rect 301890 734 302734 856
rect 302902 734 303746 856
rect 303914 734 304758 856
rect 304926 734 305770 856
rect 305938 734 306782 856
rect 306950 734 307794 856
rect 307962 734 308806 856
rect 308974 734 309818 856
rect 309986 734 310830 856
rect 310998 734 311842 856
rect 312010 734 312854 856
rect 313022 734 313866 856
rect 314034 734 314878 856
rect 315046 734 315890 856
rect 316058 734 316902 856
rect 317070 734 317914 856
rect 318082 734 318926 856
rect 319094 734 319938 856
rect 320106 734 320950 856
rect 321118 734 321962 856
rect 322130 734 322974 856
rect 323142 734 323986 856
rect 324154 734 324998 856
rect 325166 734 326010 856
rect 326178 734 327022 856
rect 327190 734 328034 856
rect 328202 734 329046 856
rect 329214 734 330058 856
rect 330226 734 331070 856
rect 331238 734 332082 856
rect 332250 734 333094 856
rect 333262 734 334106 856
rect 334274 734 335118 856
rect 335286 734 336130 856
rect 336298 734 337142 856
rect 337310 734 338154 856
rect 338322 734 339166 856
rect 339334 734 340178 856
rect 340346 734 341190 856
rect 341358 734 342202 856
rect 342370 734 343214 856
rect 343382 734 344226 856
rect 344394 734 345238 856
rect 345406 734 346250 856
rect 346418 734 347262 856
rect 347430 734 348274 856
rect 348442 734 349286 856
rect 349454 734 350298 856
rect 350466 734 351310 856
rect 351478 734 352322 856
rect 352490 734 353334 856
rect 353502 734 354346 856
rect 354514 734 355358 856
rect 355526 734 356370 856
rect 356538 734 357382 856
rect 357550 734 358394 856
rect 358562 734 359406 856
rect 359574 734 360418 856
rect 360586 734 361430 856
rect 361598 734 362442 856
rect 362610 734 363454 856
rect 363622 734 364466 856
rect 364634 734 365478 856
rect 365646 734 366490 856
rect 366658 734 367502 856
rect 367670 734 368514 856
rect 368682 734 369526 856
rect 369694 734 370538 856
rect 370706 734 371550 856
rect 371718 734 372562 856
rect 372730 734 373574 856
rect 373742 734 374586 856
rect 374754 734 375598 856
rect 375766 734 376610 856
rect 376778 734 377622 856
rect 377790 734 378634 856
rect 378802 734 379646 856
rect 379814 734 380658 856
rect 380826 734 381670 856
rect 381838 734 382682 856
rect 382850 734 383694 856
rect 383862 734 384706 856
rect 384874 734 385718 856
rect 385886 734 386730 856
rect 386898 734 387742 856
rect 387910 734 388754 856
rect 388922 734 389766 856
rect 389934 734 390778 856
rect 390946 734 391790 856
rect 391958 734 392802 856
rect 392970 734 393814 856
rect 393982 734 394826 856
rect 394994 734 395838 856
rect 396006 734 396850 856
rect 397018 734 397862 856
rect 398030 734 398874 856
rect 399042 734 399886 856
rect 400054 734 400898 856
rect 401066 734 401910 856
rect 402078 734 402922 856
rect 403090 734 403934 856
rect 404102 734 404946 856
rect 405114 734 405958 856
rect 406126 734 406970 856
rect 407138 734 407982 856
rect 408150 734 408994 856
rect 409162 734 410006 856
rect 410174 734 411018 856
rect 411186 734 412030 856
rect 412198 734 413042 856
rect 413210 734 414054 856
rect 414222 734 415066 856
rect 415234 734 416078 856
rect 416246 734 417090 856
rect 417258 734 418102 856
rect 418270 734 419114 856
rect 419282 734 420126 856
rect 420294 734 421138 856
rect 421306 734 422150 856
rect 422318 734 423162 856
rect 423330 734 424174 856
rect 424342 734 425186 856
rect 425354 734 426198 856
rect 426366 734 427210 856
rect 427378 734 428222 856
rect 428390 734 429234 856
rect 429402 734 430246 856
rect 430414 734 431258 856
rect 431426 734 432270 856
rect 432438 734 433282 856
rect 433450 734 434294 856
rect 434462 734 435306 856
rect 435474 734 436318 856
rect 436486 734 437330 856
rect 437498 734 438342 856
rect 438510 734 439354 856
rect 439522 734 440366 856
rect 440534 734 441378 856
rect 441546 734 442390 856
rect 442558 734 443402 856
rect 443570 734 444414 856
rect 444582 734 445426 856
rect 445594 734 446438 856
rect 446606 734 447450 856
rect 447618 734 448462 856
rect 448630 734 449474 856
rect 449642 734 450486 856
rect 450654 734 451498 856
rect 451666 734 452510 856
rect 452678 734 453522 856
rect 453690 734 454534 856
rect 454702 734 455546 856
rect 455714 734 456558 856
rect 456726 734 457570 856
rect 457738 734 458582 856
rect 458750 734 459594 856
rect 459762 734 460606 856
rect 460774 734 461618 856
rect 461786 734 462630 856
rect 462798 734 463642 856
rect 463810 734 464654 856
rect 464822 734 465666 856
rect 465834 734 466678 856
rect 466846 734 467690 856
rect 467858 734 468702 856
rect 468870 734 469714 856
rect 469882 734 470726 856
rect 470894 734 471738 856
rect 471906 734 472750 856
rect 472918 734 473762 856
rect 473930 734 474774 856
rect 474942 734 475786 856
rect 475954 734 476798 856
rect 476966 734 477810 856
rect 477978 734 478822 856
rect 478990 734 479834 856
rect 480002 734 480846 856
rect 481014 734 481858 856
rect 482026 734 482870 856
rect 483038 734 483882 856
rect 484050 734 484894 856
rect 485062 734 485906 856
rect 486074 734 486918 856
rect 487086 734 487930 856
rect 488098 734 488942 856
rect 489110 734 489954 856
rect 490122 734 490966 856
rect 491134 734 491978 856
rect 492146 734 492990 856
rect 493158 734 494002 856
rect 494170 734 495014 856
rect 495182 734 496026 856
rect 496194 734 497038 856
rect 497206 734 498050 856
rect 498218 734 499062 856
rect 499230 734 500074 856
rect 500242 734 501086 856
rect 501254 734 502098 856
rect 502266 734 503110 856
rect 503278 734 504122 856
rect 504290 734 505134 856
rect 505302 734 506146 856
rect 506314 734 507158 856
rect 507326 734 508170 856
rect 508338 734 509182 856
rect 509350 734 510194 856
rect 510362 734 511206 856
rect 511374 734 512218 856
rect 512386 734 513230 856
rect 513398 734 514242 856
rect 514410 734 515254 856
rect 515422 734 516266 856
rect 516434 734 517278 856
rect 517446 734 518290 856
rect 518458 734 519302 856
rect 519470 734 539010 856
<< metal3 >>
rect 0 294856 800 294976
rect 539200 293496 540000 293616
rect 0 287784 800 287904
rect 539200 286968 540000 287088
rect 0 280712 800 280832
rect 539200 280440 540000 280560
rect 539200 273912 540000 274032
rect 0 273640 800 273760
rect 539200 267384 540000 267504
rect 0 266568 800 266688
rect 539200 260856 540000 260976
rect 0 259496 800 259616
rect 539200 254328 540000 254448
rect 0 252424 800 252544
rect 539200 247800 540000 247920
rect 0 245352 800 245472
rect 539200 241272 540000 241392
rect 0 238280 800 238400
rect 539200 234744 540000 234864
rect 0 231208 800 231328
rect 539200 228216 540000 228336
rect 0 224136 800 224256
rect 539200 221688 540000 221808
rect 0 217064 800 217184
rect 539200 215160 540000 215280
rect 0 209992 800 210112
rect 539200 208632 540000 208752
rect 0 202920 800 203040
rect 539200 202104 540000 202224
rect 0 195848 800 195968
rect 539200 195576 540000 195696
rect 539200 189048 540000 189168
rect 0 188776 800 188896
rect 539200 182520 540000 182640
rect 0 181704 800 181824
rect 539200 175992 540000 176112
rect 0 174632 800 174752
rect 539200 169464 540000 169584
rect 0 167560 800 167680
rect 539200 162936 540000 163056
rect 0 160488 800 160608
rect 539200 156408 540000 156528
rect 0 153416 800 153536
rect 539200 149880 540000 150000
rect 0 146344 800 146464
rect 539200 143352 540000 143472
rect 0 139272 800 139392
rect 539200 136824 540000 136944
rect 0 132200 800 132320
rect 539200 130296 540000 130416
rect 0 125128 800 125248
rect 539200 123768 540000 123888
rect 0 118056 800 118176
rect 539200 117240 540000 117360
rect 0 110984 800 111104
rect 539200 110712 540000 110832
rect 539200 104184 540000 104304
rect 0 103912 800 104032
rect 539200 97656 540000 97776
rect 0 96840 800 96960
rect 539200 91128 540000 91248
rect 0 89768 800 89888
rect 539200 84600 540000 84720
rect 0 82696 800 82816
rect 539200 78072 540000 78192
rect 0 75624 800 75744
rect 539200 71544 540000 71664
rect 0 68552 800 68672
rect 539200 65016 540000 65136
rect 0 61480 800 61600
rect 539200 58488 540000 58608
rect 0 54408 800 54528
rect 539200 51960 540000 52080
rect 0 47336 800 47456
rect 539200 45432 540000 45552
rect 0 40264 800 40384
rect 539200 38904 540000 39024
rect 0 33192 800 33312
rect 539200 32376 540000 32496
rect 0 26120 800 26240
rect 539200 25848 540000 25968
rect 539200 19320 540000 19440
rect 0 19048 800 19168
rect 539200 12792 540000 12912
rect 0 11976 800 12096
rect 539200 6264 540000 6384
rect 0 4904 800 5024
<< obsm3 >>
rect 798 295056 539200 297601
rect 880 294776 539200 295056
rect 798 293696 539200 294776
rect 798 293416 539120 293696
rect 798 287984 539200 293416
rect 880 287704 539200 287984
rect 798 287168 539200 287704
rect 798 286888 539120 287168
rect 798 280912 539200 286888
rect 880 280640 539200 280912
rect 880 280632 539120 280640
rect 798 280360 539120 280632
rect 798 274112 539200 280360
rect 798 273840 539120 274112
rect 880 273832 539120 273840
rect 880 273560 539200 273832
rect 798 267584 539200 273560
rect 798 267304 539120 267584
rect 798 266768 539200 267304
rect 880 266488 539200 266768
rect 798 261056 539200 266488
rect 798 260776 539120 261056
rect 798 259696 539200 260776
rect 880 259416 539200 259696
rect 798 254528 539200 259416
rect 798 254248 539120 254528
rect 798 252624 539200 254248
rect 880 252344 539200 252624
rect 798 248000 539200 252344
rect 798 247720 539120 248000
rect 798 245552 539200 247720
rect 880 245272 539200 245552
rect 798 241472 539200 245272
rect 798 241192 539120 241472
rect 798 238480 539200 241192
rect 880 238200 539200 238480
rect 798 234944 539200 238200
rect 798 234664 539120 234944
rect 798 231408 539200 234664
rect 880 231128 539200 231408
rect 798 228416 539200 231128
rect 798 228136 539120 228416
rect 798 224336 539200 228136
rect 880 224056 539200 224336
rect 798 221888 539200 224056
rect 798 221608 539120 221888
rect 798 217264 539200 221608
rect 880 216984 539200 217264
rect 798 215360 539200 216984
rect 798 215080 539120 215360
rect 798 210192 539200 215080
rect 880 209912 539200 210192
rect 798 208832 539200 209912
rect 798 208552 539120 208832
rect 798 203120 539200 208552
rect 880 202840 539200 203120
rect 798 202304 539200 202840
rect 798 202024 539120 202304
rect 798 196048 539200 202024
rect 880 195776 539200 196048
rect 880 195768 539120 195776
rect 798 195496 539120 195768
rect 798 189248 539200 195496
rect 798 188976 539120 189248
rect 880 188968 539120 188976
rect 880 188696 539200 188968
rect 798 182720 539200 188696
rect 798 182440 539120 182720
rect 798 181904 539200 182440
rect 880 181624 539200 181904
rect 798 176192 539200 181624
rect 798 175912 539120 176192
rect 798 174832 539200 175912
rect 880 174552 539200 174832
rect 798 169664 539200 174552
rect 798 169384 539120 169664
rect 798 167760 539200 169384
rect 880 167480 539200 167760
rect 798 163136 539200 167480
rect 798 162856 539120 163136
rect 798 160688 539200 162856
rect 880 160408 539200 160688
rect 798 156608 539200 160408
rect 798 156328 539120 156608
rect 798 153616 539200 156328
rect 880 153336 539200 153616
rect 798 150080 539200 153336
rect 798 149800 539120 150080
rect 798 146544 539200 149800
rect 880 146264 539200 146544
rect 798 143552 539200 146264
rect 798 143272 539120 143552
rect 798 139472 539200 143272
rect 880 139192 539200 139472
rect 798 137024 539200 139192
rect 798 136744 539120 137024
rect 798 132400 539200 136744
rect 880 132120 539200 132400
rect 798 130496 539200 132120
rect 798 130216 539120 130496
rect 798 125328 539200 130216
rect 880 125048 539200 125328
rect 798 123968 539200 125048
rect 798 123688 539120 123968
rect 798 118256 539200 123688
rect 880 117976 539200 118256
rect 798 117440 539200 117976
rect 798 117160 539120 117440
rect 798 111184 539200 117160
rect 880 110912 539200 111184
rect 880 110904 539120 110912
rect 798 110632 539120 110904
rect 798 104384 539200 110632
rect 798 104112 539120 104384
rect 880 104104 539120 104112
rect 880 103832 539200 104104
rect 798 97856 539200 103832
rect 798 97576 539120 97856
rect 798 97040 539200 97576
rect 880 96760 539200 97040
rect 798 91328 539200 96760
rect 798 91048 539120 91328
rect 798 89968 539200 91048
rect 880 89688 539200 89968
rect 798 84800 539200 89688
rect 798 84520 539120 84800
rect 798 82896 539200 84520
rect 880 82616 539200 82896
rect 798 78272 539200 82616
rect 798 77992 539120 78272
rect 798 75824 539200 77992
rect 880 75544 539200 75824
rect 798 71744 539200 75544
rect 798 71464 539120 71744
rect 798 68752 539200 71464
rect 880 68472 539200 68752
rect 798 65216 539200 68472
rect 798 64936 539120 65216
rect 798 61680 539200 64936
rect 880 61400 539200 61680
rect 798 58688 539200 61400
rect 798 58408 539120 58688
rect 798 54608 539200 58408
rect 880 54328 539200 54608
rect 798 52160 539200 54328
rect 798 51880 539120 52160
rect 798 47536 539200 51880
rect 880 47256 539200 47536
rect 798 45632 539200 47256
rect 798 45352 539120 45632
rect 798 40464 539200 45352
rect 880 40184 539200 40464
rect 798 39104 539200 40184
rect 798 38824 539120 39104
rect 798 33392 539200 38824
rect 880 33112 539200 33392
rect 798 32576 539200 33112
rect 798 32296 539120 32576
rect 798 26320 539200 32296
rect 880 26048 539200 26320
rect 880 26040 539120 26048
rect 798 25768 539120 26040
rect 798 19520 539200 25768
rect 798 19248 539120 19520
rect 880 19240 539120 19248
rect 880 18968 539200 19240
rect 798 12992 539200 18968
rect 798 12712 539120 12992
rect 798 12176 539200 12712
rect 880 11896 539200 12176
rect 798 6464 539200 11896
rect 798 6184 539120 6464
rect 798 5104 539200 6184
rect 880 4824 539200 5104
rect 798 1259 539200 4824
<< metal4 >>
rect 4208 2128 4528 297616
rect 19568 2128 19888 297616
rect 34928 2128 35248 297616
rect 50288 2128 50608 297616
rect 65648 2128 65968 297616
rect 81008 2128 81328 297616
rect 96368 2128 96688 297616
rect 111728 2128 112048 297616
rect 127088 2128 127408 297616
rect 142448 2128 142768 297616
rect 157808 2128 158128 297616
rect 173168 2128 173488 297616
rect 188528 2128 188848 297616
rect 203888 2128 204208 297616
rect 219248 2128 219568 297616
rect 234608 2128 234928 297616
rect 249968 2128 250288 297616
rect 265328 2128 265648 297616
rect 280688 2128 281008 297616
rect 296048 2128 296368 297616
rect 311408 2128 311728 297616
rect 326768 2128 327088 297616
rect 342128 2128 342448 297616
rect 357488 2128 357808 297616
rect 372848 2128 373168 297616
rect 388208 2128 388528 297616
rect 403568 2128 403888 297616
rect 418928 2128 419248 297616
rect 434288 2128 434608 297616
rect 449648 2128 449968 297616
rect 465008 2128 465328 297616
rect 480368 2128 480688 297616
rect 495728 2128 496048 297616
rect 511088 2128 511408 297616
rect 526448 2128 526768 297616
<< obsm4 >>
rect 308995 38931 311328 79389
rect 311808 38931 326688 79389
rect 327168 38931 342048 79389
rect 342528 38931 357408 79389
rect 357888 38931 372768 79389
rect 373248 38931 388128 79389
rect 388608 38931 403488 79389
rect 403968 38931 415229 79389
<< labels >>
rlabel metal3 s 539200 6264 540000 6384 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 539200 202104 540000 202224 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 539200 221688 540000 221808 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 539200 241272 540000 241392 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 539200 260856 540000 260976 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 539200 280440 540000 280560 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 529478 299200 529534 300000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 469586 299200 469642 300000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 409694 299200 409750 300000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 349802 299200 349858 300000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 289910 299200 289966 300000 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 539200 25848 540000 25968 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 230018 299200 230074 300000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 170126 299200 170182 300000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 110234 299200 110290 300000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 50342 299200 50398 300000 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s 0 294856 800 294976 6 io_in[24]
port 17 nsew signal input
rlabel metal3 s 0 273640 800 273760 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 0 252424 800 252544 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 0 231208 800 231328 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 0 209992 800 210112 6 io_in[28]
port 21 nsew signal input
rlabel metal3 s 0 188776 800 188896 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 539200 45432 540000 45552 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s 0 167560 800 167680 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 0 146344 800 146464 6 io_in[31]
port 25 nsew signal input
rlabel metal3 s 0 125128 800 125248 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 0 103912 800 104032 6 io_in[33]
port 27 nsew signal input
rlabel metal3 s 0 82696 800 82816 6 io_in[34]
port 28 nsew signal input
rlabel metal3 s 0 61480 800 61600 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 0 40264 800 40384 6 io_in[36]
port 30 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 539200 65016 540000 65136 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 539200 84600 540000 84720 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 539200 104184 540000 104304 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 539200 123768 540000 123888 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 539200 143352 540000 143472 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 539200 162936 540000 163056 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 539200 182520 540000 182640 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 539200 19320 540000 19440 6 io_oeb[0]
port 39 nsew signal output
rlabel metal3 s 539200 215160 540000 215280 6 io_oeb[10]
port 40 nsew signal output
rlabel metal3 s 539200 234744 540000 234864 6 io_oeb[11]
port 41 nsew signal output
rlabel metal3 s 539200 254328 540000 254448 6 io_oeb[12]
port 42 nsew signal output
rlabel metal3 s 539200 273912 540000 274032 6 io_oeb[13]
port 43 nsew signal output
rlabel metal3 s 539200 293496 540000 293616 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 489550 299200 489606 300000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 429658 299200 429714 300000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 369766 299200 369822 300000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 309874 299200 309930 300000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 249982 299200 250038 300000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal3 s 539200 38904 540000 39024 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 190090 299200 190146 300000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 130198 299200 130254 300000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 70306 299200 70362 300000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 10414 299200 10470 300000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s 0 280712 800 280832 6 io_oeb[24]
port 55 nsew signal output
rlabel metal3 s 0 259496 800 259616 6 io_oeb[25]
port 56 nsew signal output
rlabel metal3 s 0 238280 800 238400 6 io_oeb[26]
port 57 nsew signal output
rlabel metal3 s 0 217064 800 217184 6 io_oeb[27]
port 58 nsew signal output
rlabel metal3 s 0 195848 800 195968 6 io_oeb[28]
port 59 nsew signal output
rlabel metal3 s 0 174632 800 174752 6 io_oeb[29]
port 60 nsew signal output
rlabel metal3 s 539200 58488 540000 58608 6 io_oeb[2]
port 61 nsew signal output
rlabel metal3 s 0 153416 800 153536 6 io_oeb[30]
port 62 nsew signal output
rlabel metal3 s 0 132200 800 132320 6 io_oeb[31]
port 63 nsew signal output
rlabel metal3 s 0 110984 800 111104 6 io_oeb[32]
port 64 nsew signal output
rlabel metal3 s 0 89768 800 89888 6 io_oeb[33]
port 65 nsew signal output
rlabel metal3 s 0 68552 800 68672 6 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s 0 47336 800 47456 6 io_oeb[35]
port 67 nsew signal output
rlabel metal3 s 0 26120 800 26240 6 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s 0 4904 800 5024 6 io_oeb[37]
port 69 nsew signal output
rlabel metal3 s 539200 78072 540000 78192 6 io_oeb[3]
port 70 nsew signal output
rlabel metal3 s 539200 97656 540000 97776 6 io_oeb[4]
port 71 nsew signal output
rlabel metal3 s 539200 117240 540000 117360 6 io_oeb[5]
port 72 nsew signal output
rlabel metal3 s 539200 136824 540000 136944 6 io_oeb[6]
port 73 nsew signal output
rlabel metal3 s 539200 156408 540000 156528 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 539200 175992 540000 176112 6 io_oeb[8]
port 75 nsew signal output
rlabel metal3 s 539200 195576 540000 195696 6 io_oeb[9]
port 76 nsew signal output
rlabel metal3 s 539200 12792 540000 12912 6 io_out[0]
port 77 nsew signal output
rlabel metal3 s 539200 208632 540000 208752 6 io_out[10]
port 78 nsew signal output
rlabel metal3 s 539200 228216 540000 228336 6 io_out[11]
port 79 nsew signal output
rlabel metal3 s 539200 247800 540000 247920 6 io_out[12]
port 80 nsew signal output
rlabel metal3 s 539200 267384 540000 267504 6 io_out[13]
port 81 nsew signal output
rlabel metal3 s 539200 286968 540000 287088 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 509514 299200 509570 300000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 449622 299200 449678 300000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 389730 299200 389786 300000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 329838 299200 329894 300000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 269946 299200 270002 300000 6 io_out[19]
port 87 nsew signal output
rlabel metal3 s 539200 32376 540000 32496 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 210054 299200 210110 300000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 150162 299200 150218 300000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 90270 299200 90326 300000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 30378 299200 30434 300000 6 io_out[23]
port 92 nsew signal output
rlabel metal3 s 0 287784 800 287904 6 io_out[24]
port 93 nsew signal output
rlabel metal3 s 0 266568 800 266688 6 io_out[25]
port 94 nsew signal output
rlabel metal3 s 0 245352 800 245472 6 io_out[26]
port 95 nsew signal output
rlabel metal3 s 0 224136 800 224256 6 io_out[27]
port 96 nsew signal output
rlabel metal3 s 0 202920 800 203040 6 io_out[28]
port 97 nsew signal output
rlabel metal3 s 0 181704 800 181824 6 io_out[29]
port 98 nsew signal output
rlabel metal3 s 539200 51960 540000 52080 6 io_out[2]
port 99 nsew signal output
rlabel metal3 s 0 160488 800 160608 6 io_out[30]
port 100 nsew signal output
rlabel metal3 s 0 139272 800 139392 6 io_out[31]
port 101 nsew signal output
rlabel metal3 s 0 118056 800 118176 6 io_out[32]
port 102 nsew signal output
rlabel metal3 s 0 96840 800 96960 6 io_out[33]
port 103 nsew signal output
rlabel metal3 s 0 75624 800 75744 6 io_out[34]
port 104 nsew signal output
rlabel metal3 s 0 54408 800 54528 6 io_out[35]
port 105 nsew signal output
rlabel metal3 s 0 33192 800 33312 6 io_out[36]
port 106 nsew signal output
rlabel metal3 s 0 11976 800 12096 6 io_out[37]
port 107 nsew signal output
rlabel metal3 s 539200 71544 540000 71664 6 io_out[3]
port 108 nsew signal output
rlabel metal3 s 539200 91128 540000 91248 6 io_out[4]
port 109 nsew signal output
rlabel metal3 s 539200 110712 540000 110832 6 io_out[5]
port 110 nsew signal output
rlabel metal3 s 539200 130296 540000 130416 6 io_out[6]
port 111 nsew signal output
rlabel metal3 s 539200 149880 540000 150000 6 io_out[7]
port 112 nsew signal output
rlabel metal3 s 539200 169464 540000 169584 6 io_out[8]
port 113 nsew signal output
rlabel metal3 s 539200 189048 540000 189168 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 516322 0 516378 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 517334 0 517390 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 518346 0 518402 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 127714 0 127770 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 431314 0 431370 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 434350 0 434406 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 437386 0 437442 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 440422 0 440478 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 443458 0 443514 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 446494 0 446550 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 449530 0 449586 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 452566 0 452622 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 455602 0 455658 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 458638 0 458694 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 158074 0 158130 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 461674 0 461730 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 464710 0 464766 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 467746 0 467802 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 470782 0 470838 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 473818 0 473874 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 476854 0 476910 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 479890 0 479946 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 482926 0 482982 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 485962 0 486018 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 488998 0 489054 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 161110 0 161166 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 492034 0 492090 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 495070 0 495126 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 498106 0 498162 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 501142 0 501198 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 504178 0 504234 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 507214 0 507270 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 510250 0 510306 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 513286 0 513342 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 164146 0 164202 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 167182 0 167238 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 170218 0 170274 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 173254 0 173310 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 176290 0 176346 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 179326 0 179382 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 182362 0 182418 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 185398 0 185454 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 130750 0 130806 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 188434 0 188490 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 191470 0 191526 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 194506 0 194562 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 197542 0 197598 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 200578 0 200634 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 203614 0 203670 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 206650 0 206706 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 209686 0 209742 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 212722 0 212778 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 215758 0 215814 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 133786 0 133842 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 218794 0 218850 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 221830 0 221886 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 224866 0 224922 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 227902 0 227958 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 230938 0 230994 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 233974 0 234030 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 237010 0 237066 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 240046 0 240102 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 243082 0 243138 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 246118 0 246174 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 136822 0 136878 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 249154 0 249210 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 252190 0 252246 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 255226 0 255282 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 258262 0 258318 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 261298 0 261354 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 264334 0 264390 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 267370 0 267426 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 270406 0 270462 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 273442 0 273498 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 276478 0 276534 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 139858 0 139914 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 279514 0 279570 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 282550 0 282606 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 285586 0 285642 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 288622 0 288678 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 291658 0 291714 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 294694 0 294750 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 297730 0 297786 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 300766 0 300822 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 303802 0 303858 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 306838 0 306894 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 142894 0 142950 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 309874 0 309930 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 312910 0 312966 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 315946 0 316002 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 318982 0 319038 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 322018 0 322074 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 325054 0 325110 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 328090 0 328146 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 331126 0 331182 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 334162 0 334218 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 337198 0 337254 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 145930 0 145986 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 340234 0 340290 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 343270 0 343326 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 346306 0 346362 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 349342 0 349398 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 352378 0 352434 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 355414 0 355470 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 358450 0 358506 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 361486 0 361542 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 364522 0 364578 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 367558 0 367614 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 148966 0 149022 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 370594 0 370650 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 373630 0 373686 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 376666 0 376722 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 379702 0 379758 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 382738 0 382794 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 385774 0 385830 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 388810 0 388866 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 391846 0 391902 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 394882 0 394938 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 397918 0 397974 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 152002 0 152058 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 400954 0 401010 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 403990 0 404046 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 407026 0 407082 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 410062 0 410118 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 413098 0 413154 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 416134 0 416190 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 419170 0 419226 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 422206 0 422262 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 425242 0 425298 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 428278 0 428334 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 155038 0 155094 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 128726 0 128782 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 432326 0 432382 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 435362 0 435418 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 438398 0 438454 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 441434 0 441490 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 444470 0 444526 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 447506 0 447562 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 450542 0 450598 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 453578 0 453634 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 456614 0 456670 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 459650 0 459706 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 159086 0 159142 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 462686 0 462742 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 465722 0 465778 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 468758 0 468814 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 471794 0 471850 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 474830 0 474886 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 477866 0 477922 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 480902 0 480958 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 483938 0 483994 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 486974 0 487030 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 490010 0 490066 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 162122 0 162178 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 493046 0 493102 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 496082 0 496138 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 499118 0 499174 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 502154 0 502210 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 505190 0 505246 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 508226 0 508282 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 511262 0 511318 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 514298 0 514354 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 165158 0 165214 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 168194 0 168250 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 171230 0 171286 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 174266 0 174322 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 177302 0 177358 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 180338 0 180394 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 183374 0 183430 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 186410 0 186466 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 131762 0 131818 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 189446 0 189502 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 192482 0 192538 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 195518 0 195574 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 198554 0 198610 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 201590 0 201646 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 204626 0 204682 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 207662 0 207718 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 210698 0 210754 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 213734 0 213790 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 216770 0 216826 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 134798 0 134854 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 219806 0 219862 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 222842 0 222898 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 225878 0 225934 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 228914 0 228970 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 231950 0 232006 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 234986 0 235042 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 238022 0 238078 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 241058 0 241114 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 244094 0 244150 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 247130 0 247186 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 137834 0 137890 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 250166 0 250222 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 253202 0 253258 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 256238 0 256294 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 259274 0 259330 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 262310 0 262366 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 265346 0 265402 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 268382 0 268438 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 271418 0 271474 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 274454 0 274510 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 277490 0 277546 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 140870 0 140926 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 280526 0 280582 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 283562 0 283618 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 286598 0 286654 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 289634 0 289690 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 292670 0 292726 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 295706 0 295762 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 298742 0 298798 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 301778 0 301834 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 304814 0 304870 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 307850 0 307906 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 143906 0 143962 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 310886 0 310942 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 313922 0 313978 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 316958 0 317014 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 319994 0 320050 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 323030 0 323086 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 326066 0 326122 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 329102 0 329158 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 332138 0 332194 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 335174 0 335230 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 338210 0 338266 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 146942 0 146998 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 341246 0 341302 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 344282 0 344338 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 347318 0 347374 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 350354 0 350410 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 353390 0 353446 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 356426 0 356482 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 359462 0 359518 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 362498 0 362554 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 365534 0 365590 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 368570 0 368626 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 149978 0 150034 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 371606 0 371662 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 374642 0 374698 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 377678 0 377734 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 380714 0 380770 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 383750 0 383806 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 386786 0 386842 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 389822 0 389878 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 392858 0 392914 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 395894 0 395950 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 398930 0 398986 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 153014 0 153070 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 401966 0 402022 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 405002 0 405058 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 408038 0 408094 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 411074 0 411130 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 414110 0 414166 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 417146 0 417202 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 420182 0 420238 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 423218 0 423274 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 426254 0 426310 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 429290 0 429346 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 156050 0 156106 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 129738 0 129794 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 433338 0 433394 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 436374 0 436430 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 439410 0 439466 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 442446 0 442502 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 445482 0 445538 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 448518 0 448574 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 451554 0 451610 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 454590 0 454646 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 457626 0 457682 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 460662 0 460718 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 160098 0 160154 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 463698 0 463754 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 466734 0 466790 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 469770 0 469826 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 472806 0 472862 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 475842 0 475898 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 478878 0 478934 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 481914 0 481970 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 484950 0 485006 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 487986 0 488042 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 491022 0 491078 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 163134 0 163190 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 494058 0 494114 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 497094 0 497150 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 500130 0 500186 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 503166 0 503222 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 506202 0 506258 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 509238 0 509294 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 512274 0 512330 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 515310 0 515366 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 166170 0 166226 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 169206 0 169262 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 172242 0 172298 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 175278 0 175334 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 178314 0 178370 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 181350 0 181406 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 184386 0 184442 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 187422 0 187478 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 132774 0 132830 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 190458 0 190514 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 193494 0 193550 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 196530 0 196586 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 199566 0 199622 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 202602 0 202658 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 205638 0 205694 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 208674 0 208730 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 211710 0 211766 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 214746 0 214802 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 217782 0 217838 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 135810 0 135866 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 220818 0 220874 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 223854 0 223910 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 226890 0 226946 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 229926 0 229982 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 232962 0 233018 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 235998 0 236054 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 239034 0 239090 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 242070 0 242126 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 245106 0 245162 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 248142 0 248198 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 138846 0 138902 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 251178 0 251234 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 254214 0 254270 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 257250 0 257306 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 260286 0 260342 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 263322 0 263378 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 266358 0 266414 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 269394 0 269450 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 272430 0 272486 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 275466 0 275522 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 278502 0 278558 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 141882 0 141938 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 281538 0 281594 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 284574 0 284630 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 287610 0 287666 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 290646 0 290702 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 293682 0 293738 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 296718 0 296774 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 299754 0 299810 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 302790 0 302846 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 305826 0 305882 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 308862 0 308918 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 144918 0 144974 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 311898 0 311954 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 314934 0 314990 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 317970 0 318026 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 321006 0 321062 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 324042 0 324098 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 327078 0 327134 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 330114 0 330170 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 333150 0 333206 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 336186 0 336242 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 339222 0 339278 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 147954 0 148010 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 342258 0 342314 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 345294 0 345350 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 348330 0 348386 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 351366 0 351422 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 354402 0 354458 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 357438 0 357494 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 360474 0 360530 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 363510 0 363566 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 366546 0 366602 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 369582 0 369638 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 150990 0 151046 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 372618 0 372674 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 375654 0 375710 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 378690 0 378746 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 381726 0 381782 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 384762 0 384818 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 387798 0 387854 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 390834 0 390890 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 393870 0 393926 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 396906 0 396962 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 399942 0 399998 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 154026 0 154082 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 402978 0 403034 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 406014 0 406070 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 409050 0 409106 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 412086 0 412142 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 415122 0 415178 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 418158 0 418214 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 421194 0 421250 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 424230 0 424286 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 427266 0 427322 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 430302 0 430358 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 157062 0 157118 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal2 s 519358 0 519414 800 6 user_clock2
port 502 nsew signal input
rlabel metal4 s 4208 2128 4528 297616 6 vccd1
port 503 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 297616 6 vccd1
port 503 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 297616 6 vccd1
port 503 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 297616 6 vccd1
port 503 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 297616 6 vccd1
port 503 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 297616 6 vccd1
port 503 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 297616 6 vccd1
port 503 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 297616 6 vccd1
port 503 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 297616 6 vccd1
port 503 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 297616 6 vccd1
port 503 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 297616 6 vccd1
port 503 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 297616 6 vccd1
port 503 nsew power bidirectional
rlabel metal4 s 372848 2128 373168 297616 6 vccd1
port 503 nsew power bidirectional
rlabel metal4 s 403568 2128 403888 297616 6 vccd1
port 503 nsew power bidirectional
rlabel metal4 s 434288 2128 434608 297616 6 vccd1
port 503 nsew power bidirectional
rlabel metal4 s 465008 2128 465328 297616 6 vccd1
port 503 nsew power bidirectional
rlabel metal4 s 495728 2128 496048 297616 6 vccd1
port 503 nsew power bidirectional
rlabel metal4 s 526448 2128 526768 297616 6 vccd1
port 503 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 297616 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 297616 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 297616 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 297616 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 297616 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 297616 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 297616 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 297616 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 297616 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 297616 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 297616 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 357488 2128 357808 297616 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 388208 2128 388528 297616 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 418928 2128 419248 297616 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 449648 2128 449968 297616 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 480368 2128 480688 297616 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 511088 2128 511408 297616 6 vssd1
port 504 nsew ground bidirectional
rlabel metal2 s 20442 0 20498 800 6 wb_clk_i
port 505 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 wb_rst_i
port 506 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 wbs_ack_o
port 507 nsew signal output
rlabel metal2 s 26514 0 26570 800 6 wbs_adr_i[0]
port 508 nsew signal input
rlabel metal2 s 60922 0 60978 800 6 wbs_adr_i[10]
port 509 nsew signal input
rlabel metal2 s 63958 0 64014 800 6 wbs_adr_i[11]
port 510 nsew signal input
rlabel metal2 s 66994 0 67050 800 6 wbs_adr_i[12]
port 511 nsew signal input
rlabel metal2 s 70030 0 70086 800 6 wbs_adr_i[13]
port 512 nsew signal input
rlabel metal2 s 73066 0 73122 800 6 wbs_adr_i[14]
port 513 nsew signal input
rlabel metal2 s 76102 0 76158 800 6 wbs_adr_i[15]
port 514 nsew signal input
rlabel metal2 s 79138 0 79194 800 6 wbs_adr_i[16]
port 515 nsew signal input
rlabel metal2 s 82174 0 82230 800 6 wbs_adr_i[17]
port 516 nsew signal input
rlabel metal2 s 85210 0 85266 800 6 wbs_adr_i[18]
port 517 nsew signal input
rlabel metal2 s 88246 0 88302 800 6 wbs_adr_i[19]
port 518 nsew signal input
rlabel metal2 s 30562 0 30618 800 6 wbs_adr_i[1]
port 519 nsew signal input
rlabel metal2 s 91282 0 91338 800 6 wbs_adr_i[20]
port 520 nsew signal input
rlabel metal2 s 94318 0 94374 800 6 wbs_adr_i[21]
port 521 nsew signal input
rlabel metal2 s 97354 0 97410 800 6 wbs_adr_i[22]
port 522 nsew signal input
rlabel metal2 s 100390 0 100446 800 6 wbs_adr_i[23]
port 523 nsew signal input
rlabel metal2 s 103426 0 103482 800 6 wbs_adr_i[24]
port 524 nsew signal input
rlabel metal2 s 106462 0 106518 800 6 wbs_adr_i[25]
port 525 nsew signal input
rlabel metal2 s 109498 0 109554 800 6 wbs_adr_i[26]
port 526 nsew signal input
rlabel metal2 s 112534 0 112590 800 6 wbs_adr_i[27]
port 527 nsew signal input
rlabel metal2 s 115570 0 115626 800 6 wbs_adr_i[28]
port 528 nsew signal input
rlabel metal2 s 118606 0 118662 800 6 wbs_adr_i[29]
port 529 nsew signal input
rlabel metal2 s 34610 0 34666 800 6 wbs_adr_i[2]
port 530 nsew signal input
rlabel metal2 s 121642 0 121698 800 6 wbs_adr_i[30]
port 531 nsew signal input
rlabel metal2 s 124678 0 124734 800 6 wbs_adr_i[31]
port 532 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 wbs_adr_i[3]
port 533 nsew signal input
rlabel metal2 s 42706 0 42762 800 6 wbs_adr_i[4]
port 534 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 wbs_adr_i[5]
port 535 nsew signal input
rlabel metal2 s 48778 0 48834 800 6 wbs_adr_i[6]
port 536 nsew signal input
rlabel metal2 s 51814 0 51870 800 6 wbs_adr_i[7]
port 537 nsew signal input
rlabel metal2 s 54850 0 54906 800 6 wbs_adr_i[8]
port 538 nsew signal input
rlabel metal2 s 57886 0 57942 800 6 wbs_adr_i[9]
port 539 nsew signal input
rlabel metal2 s 23478 0 23534 800 6 wbs_cyc_i
port 540 nsew signal input
rlabel metal2 s 27526 0 27582 800 6 wbs_dat_i[0]
port 541 nsew signal input
rlabel metal2 s 61934 0 61990 800 6 wbs_dat_i[10]
port 542 nsew signal input
rlabel metal2 s 64970 0 65026 800 6 wbs_dat_i[11]
port 543 nsew signal input
rlabel metal2 s 68006 0 68062 800 6 wbs_dat_i[12]
port 544 nsew signal input
rlabel metal2 s 71042 0 71098 800 6 wbs_dat_i[13]
port 545 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 wbs_dat_i[14]
port 546 nsew signal input
rlabel metal2 s 77114 0 77170 800 6 wbs_dat_i[15]
port 547 nsew signal input
rlabel metal2 s 80150 0 80206 800 6 wbs_dat_i[16]
port 548 nsew signal input
rlabel metal2 s 83186 0 83242 800 6 wbs_dat_i[17]
port 549 nsew signal input
rlabel metal2 s 86222 0 86278 800 6 wbs_dat_i[18]
port 550 nsew signal input
rlabel metal2 s 89258 0 89314 800 6 wbs_dat_i[19]
port 551 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 wbs_dat_i[1]
port 552 nsew signal input
rlabel metal2 s 92294 0 92350 800 6 wbs_dat_i[20]
port 553 nsew signal input
rlabel metal2 s 95330 0 95386 800 6 wbs_dat_i[21]
port 554 nsew signal input
rlabel metal2 s 98366 0 98422 800 6 wbs_dat_i[22]
port 555 nsew signal input
rlabel metal2 s 101402 0 101458 800 6 wbs_dat_i[23]
port 556 nsew signal input
rlabel metal2 s 104438 0 104494 800 6 wbs_dat_i[24]
port 557 nsew signal input
rlabel metal2 s 107474 0 107530 800 6 wbs_dat_i[25]
port 558 nsew signal input
rlabel metal2 s 110510 0 110566 800 6 wbs_dat_i[26]
port 559 nsew signal input
rlabel metal2 s 113546 0 113602 800 6 wbs_dat_i[27]
port 560 nsew signal input
rlabel metal2 s 116582 0 116638 800 6 wbs_dat_i[28]
port 561 nsew signal input
rlabel metal2 s 119618 0 119674 800 6 wbs_dat_i[29]
port 562 nsew signal input
rlabel metal2 s 35622 0 35678 800 6 wbs_dat_i[2]
port 563 nsew signal input
rlabel metal2 s 122654 0 122710 800 6 wbs_dat_i[30]
port 564 nsew signal input
rlabel metal2 s 125690 0 125746 800 6 wbs_dat_i[31]
port 565 nsew signal input
rlabel metal2 s 39670 0 39726 800 6 wbs_dat_i[3]
port 566 nsew signal input
rlabel metal2 s 43718 0 43774 800 6 wbs_dat_i[4]
port 567 nsew signal input
rlabel metal2 s 46754 0 46810 800 6 wbs_dat_i[5]
port 568 nsew signal input
rlabel metal2 s 49790 0 49846 800 6 wbs_dat_i[6]
port 569 nsew signal input
rlabel metal2 s 52826 0 52882 800 6 wbs_dat_i[7]
port 570 nsew signal input
rlabel metal2 s 55862 0 55918 800 6 wbs_dat_i[8]
port 571 nsew signal input
rlabel metal2 s 58898 0 58954 800 6 wbs_dat_i[9]
port 572 nsew signal input
rlabel metal2 s 28538 0 28594 800 6 wbs_dat_o[0]
port 573 nsew signal output
rlabel metal2 s 62946 0 63002 800 6 wbs_dat_o[10]
port 574 nsew signal output
rlabel metal2 s 65982 0 66038 800 6 wbs_dat_o[11]
port 575 nsew signal output
rlabel metal2 s 69018 0 69074 800 6 wbs_dat_o[12]
port 576 nsew signal output
rlabel metal2 s 72054 0 72110 800 6 wbs_dat_o[13]
port 577 nsew signal output
rlabel metal2 s 75090 0 75146 800 6 wbs_dat_o[14]
port 578 nsew signal output
rlabel metal2 s 78126 0 78182 800 6 wbs_dat_o[15]
port 579 nsew signal output
rlabel metal2 s 81162 0 81218 800 6 wbs_dat_o[16]
port 580 nsew signal output
rlabel metal2 s 84198 0 84254 800 6 wbs_dat_o[17]
port 581 nsew signal output
rlabel metal2 s 87234 0 87290 800 6 wbs_dat_o[18]
port 582 nsew signal output
rlabel metal2 s 90270 0 90326 800 6 wbs_dat_o[19]
port 583 nsew signal output
rlabel metal2 s 32586 0 32642 800 6 wbs_dat_o[1]
port 584 nsew signal output
rlabel metal2 s 93306 0 93362 800 6 wbs_dat_o[20]
port 585 nsew signal output
rlabel metal2 s 96342 0 96398 800 6 wbs_dat_o[21]
port 586 nsew signal output
rlabel metal2 s 99378 0 99434 800 6 wbs_dat_o[22]
port 587 nsew signal output
rlabel metal2 s 102414 0 102470 800 6 wbs_dat_o[23]
port 588 nsew signal output
rlabel metal2 s 105450 0 105506 800 6 wbs_dat_o[24]
port 589 nsew signal output
rlabel metal2 s 108486 0 108542 800 6 wbs_dat_o[25]
port 590 nsew signal output
rlabel metal2 s 111522 0 111578 800 6 wbs_dat_o[26]
port 591 nsew signal output
rlabel metal2 s 114558 0 114614 800 6 wbs_dat_o[27]
port 592 nsew signal output
rlabel metal2 s 117594 0 117650 800 6 wbs_dat_o[28]
port 593 nsew signal output
rlabel metal2 s 120630 0 120686 800 6 wbs_dat_o[29]
port 594 nsew signal output
rlabel metal2 s 36634 0 36690 800 6 wbs_dat_o[2]
port 595 nsew signal output
rlabel metal2 s 123666 0 123722 800 6 wbs_dat_o[30]
port 596 nsew signal output
rlabel metal2 s 126702 0 126758 800 6 wbs_dat_o[31]
port 597 nsew signal output
rlabel metal2 s 40682 0 40738 800 6 wbs_dat_o[3]
port 598 nsew signal output
rlabel metal2 s 44730 0 44786 800 6 wbs_dat_o[4]
port 599 nsew signal output
rlabel metal2 s 47766 0 47822 800 6 wbs_dat_o[5]
port 600 nsew signal output
rlabel metal2 s 50802 0 50858 800 6 wbs_dat_o[6]
port 601 nsew signal output
rlabel metal2 s 53838 0 53894 800 6 wbs_dat_o[7]
port 602 nsew signal output
rlabel metal2 s 56874 0 56930 800 6 wbs_dat_o[8]
port 603 nsew signal output
rlabel metal2 s 59910 0 59966 800 6 wbs_dat_o[9]
port 604 nsew signal output
rlabel metal2 s 29550 0 29606 800 6 wbs_sel_i[0]
port 605 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 wbs_sel_i[1]
port 606 nsew signal input
rlabel metal2 s 37646 0 37702 800 6 wbs_sel_i[2]
port 607 nsew signal input
rlabel metal2 s 41694 0 41750 800 6 wbs_sel_i[3]
port 608 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 wbs_stb_i
port 609 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 wbs_we_i
port 610 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 540000 300000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 133706762
string GDS_FILE /home/anton/projects/CUP-algofoogle/openlane/user_proj_example/runs/24_09_26_07_57/results/signoff/user_proj_example.magic.gds
string GDS_START 1177876
<< end >>

