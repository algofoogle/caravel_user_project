magic
tech sky130A
magscale 1 2
timestamp 1727137714
<< obsli1 >>
rect 1104 2159 538844 317713
<< obsm1 >>
rect 934 76 539014 317744
<< metal2 >>
rect 10414 319200 10470 320000
rect 30378 319200 30434 320000
rect 50342 319200 50398 320000
rect 70306 319200 70362 320000
rect 90270 319200 90326 320000
rect 110234 319200 110290 320000
rect 130198 319200 130254 320000
rect 150162 319200 150218 320000
rect 170126 319200 170182 320000
rect 190090 319200 190146 320000
rect 210054 319200 210110 320000
rect 230018 319200 230074 320000
rect 249982 319200 250038 320000
rect 269946 319200 270002 320000
rect 289910 319200 289966 320000
rect 309874 319200 309930 320000
rect 329838 319200 329894 320000
rect 349802 319200 349858 320000
rect 369766 319200 369822 320000
rect 389730 319200 389786 320000
rect 409694 319200 409750 320000
rect 429658 319200 429714 320000
rect 449622 319200 449678 320000
rect 469586 319200 469642 320000
rect 489550 319200 489606 320000
rect 509514 319200 509570 320000
rect 529478 319200 529534 320000
rect 20994 0 21050 800
rect 22006 0 22062 800
rect 23018 0 23074 800
rect 24030 0 24086 800
rect 25042 0 25098 800
rect 26054 0 26110 800
rect 27066 0 27122 800
rect 28078 0 28134 800
rect 29090 0 29146 800
rect 30102 0 30158 800
rect 31114 0 31170 800
rect 32126 0 32182 800
rect 33138 0 33194 800
rect 34150 0 34206 800
rect 35162 0 35218 800
rect 36174 0 36230 800
rect 37186 0 37242 800
rect 38198 0 38254 800
rect 39210 0 39266 800
rect 40222 0 40278 800
rect 41234 0 41290 800
rect 42246 0 42302 800
rect 43258 0 43314 800
rect 44270 0 44326 800
rect 45282 0 45338 800
rect 46294 0 46350 800
rect 47306 0 47362 800
rect 48318 0 48374 800
rect 49330 0 49386 800
rect 50342 0 50398 800
rect 51354 0 51410 800
rect 52366 0 52422 800
rect 53378 0 53434 800
rect 54390 0 54446 800
rect 55402 0 55458 800
rect 56414 0 56470 800
rect 57426 0 57482 800
rect 58438 0 58494 800
rect 59450 0 59506 800
rect 60462 0 60518 800
rect 61474 0 61530 800
rect 62486 0 62542 800
rect 63498 0 63554 800
rect 64510 0 64566 800
rect 65522 0 65578 800
rect 66534 0 66590 800
rect 67546 0 67602 800
rect 68558 0 68614 800
rect 69570 0 69626 800
rect 70582 0 70638 800
rect 71594 0 71650 800
rect 72606 0 72662 800
rect 73618 0 73674 800
rect 74630 0 74686 800
rect 75642 0 75698 800
rect 76654 0 76710 800
rect 77666 0 77722 800
rect 78678 0 78734 800
rect 79690 0 79746 800
rect 80702 0 80758 800
rect 81714 0 81770 800
rect 82726 0 82782 800
rect 83738 0 83794 800
rect 84750 0 84806 800
rect 85762 0 85818 800
rect 86774 0 86830 800
rect 87786 0 87842 800
rect 88798 0 88854 800
rect 89810 0 89866 800
rect 90822 0 90878 800
rect 91834 0 91890 800
rect 92846 0 92902 800
rect 93858 0 93914 800
rect 94870 0 94926 800
rect 95882 0 95938 800
rect 96894 0 96950 800
rect 97906 0 97962 800
rect 98918 0 98974 800
rect 99930 0 99986 800
rect 100942 0 100998 800
rect 101954 0 102010 800
rect 102966 0 103022 800
rect 103978 0 104034 800
rect 104990 0 105046 800
rect 106002 0 106058 800
rect 107014 0 107070 800
rect 108026 0 108082 800
rect 109038 0 109094 800
rect 110050 0 110106 800
rect 111062 0 111118 800
rect 112074 0 112130 800
rect 113086 0 113142 800
rect 114098 0 114154 800
rect 115110 0 115166 800
rect 116122 0 116178 800
rect 117134 0 117190 800
rect 118146 0 118202 800
rect 119158 0 119214 800
rect 120170 0 120226 800
rect 121182 0 121238 800
rect 122194 0 122250 800
rect 123206 0 123262 800
rect 124218 0 124274 800
rect 125230 0 125286 800
rect 126242 0 126298 800
rect 127254 0 127310 800
rect 128266 0 128322 800
rect 129278 0 129334 800
rect 130290 0 130346 800
rect 131302 0 131358 800
rect 132314 0 132370 800
rect 133326 0 133382 800
rect 134338 0 134394 800
rect 135350 0 135406 800
rect 136362 0 136418 800
rect 137374 0 137430 800
rect 138386 0 138442 800
rect 139398 0 139454 800
rect 140410 0 140466 800
rect 141422 0 141478 800
rect 142434 0 142490 800
rect 143446 0 143502 800
rect 144458 0 144514 800
rect 145470 0 145526 800
rect 146482 0 146538 800
rect 147494 0 147550 800
rect 148506 0 148562 800
rect 149518 0 149574 800
rect 150530 0 150586 800
rect 151542 0 151598 800
rect 152554 0 152610 800
rect 153566 0 153622 800
rect 154578 0 154634 800
rect 155590 0 155646 800
rect 156602 0 156658 800
rect 157614 0 157670 800
rect 158626 0 158682 800
rect 159638 0 159694 800
rect 160650 0 160706 800
rect 161662 0 161718 800
rect 162674 0 162730 800
rect 163686 0 163742 800
rect 164698 0 164754 800
rect 165710 0 165766 800
rect 166722 0 166778 800
rect 167734 0 167790 800
rect 168746 0 168802 800
rect 169758 0 169814 800
rect 170770 0 170826 800
rect 171782 0 171838 800
rect 172794 0 172850 800
rect 173806 0 173862 800
rect 174818 0 174874 800
rect 175830 0 175886 800
rect 176842 0 176898 800
rect 177854 0 177910 800
rect 178866 0 178922 800
rect 179878 0 179934 800
rect 180890 0 180946 800
rect 181902 0 181958 800
rect 182914 0 182970 800
rect 183926 0 183982 800
rect 184938 0 184994 800
rect 185950 0 186006 800
rect 186962 0 187018 800
rect 187974 0 188030 800
rect 188986 0 189042 800
rect 189998 0 190054 800
rect 191010 0 191066 800
rect 192022 0 192078 800
rect 193034 0 193090 800
rect 194046 0 194102 800
rect 195058 0 195114 800
rect 196070 0 196126 800
rect 197082 0 197138 800
rect 198094 0 198150 800
rect 199106 0 199162 800
rect 200118 0 200174 800
rect 201130 0 201186 800
rect 202142 0 202198 800
rect 203154 0 203210 800
rect 204166 0 204222 800
rect 205178 0 205234 800
rect 206190 0 206246 800
rect 207202 0 207258 800
rect 208214 0 208270 800
rect 209226 0 209282 800
rect 210238 0 210294 800
rect 211250 0 211306 800
rect 212262 0 212318 800
rect 213274 0 213330 800
rect 214286 0 214342 800
rect 215298 0 215354 800
rect 216310 0 216366 800
rect 217322 0 217378 800
rect 218334 0 218390 800
rect 219346 0 219402 800
rect 220358 0 220414 800
rect 221370 0 221426 800
rect 222382 0 222438 800
rect 223394 0 223450 800
rect 224406 0 224462 800
rect 225418 0 225474 800
rect 226430 0 226486 800
rect 227442 0 227498 800
rect 228454 0 228510 800
rect 229466 0 229522 800
rect 230478 0 230534 800
rect 231490 0 231546 800
rect 232502 0 232558 800
rect 233514 0 233570 800
rect 234526 0 234582 800
rect 235538 0 235594 800
rect 236550 0 236606 800
rect 237562 0 237618 800
rect 238574 0 238630 800
rect 239586 0 239642 800
rect 240598 0 240654 800
rect 241610 0 241666 800
rect 242622 0 242678 800
rect 243634 0 243690 800
rect 244646 0 244702 800
rect 245658 0 245714 800
rect 246670 0 246726 800
rect 247682 0 247738 800
rect 248694 0 248750 800
rect 249706 0 249762 800
rect 250718 0 250774 800
rect 251730 0 251786 800
rect 252742 0 252798 800
rect 253754 0 253810 800
rect 254766 0 254822 800
rect 255778 0 255834 800
rect 256790 0 256846 800
rect 257802 0 257858 800
rect 258814 0 258870 800
rect 259826 0 259882 800
rect 260838 0 260894 800
rect 261850 0 261906 800
rect 262862 0 262918 800
rect 263874 0 263930 800
rect 264886 0 264942 800
rect 265898 0 265954 800
rect 266910 0 266966 800
rect 267922 0 267978 800
rect 268934 0 268990 800
rect 269946 0 270002 800
rect 270958 0 271014 800
rect 271970 0 272026 800
rect 272982 0 273038 800
rect 273994 0 274050 800
rect 275006 0 275062 800
rect 276018 0 276074 800
rect 277030 0 277086 800
rect 278042 0 278098 800
rect 279054 0 279110 800
rect 280066 0 280122 800
rect 281078 0 281134 800
rect 282090 0 282146 800
rect 283102 0 283158 800
rect 284114 0 284170 800
rect 285126 0 285182 800
rect 286138 0 286194 800
rect 287150 0 287206 800
rect 288162 0 288218 800
rect 289174 0 289230 800
rect 290186 0 290242 800
rect 291198 0 291254 800
rect 292210 0 292266 800
rect 293222 0 293278 800
rect 294234 0 294290 800
rect 295246 0 295302 800
rect 296258 0 296314 800
rect 297270 0 297326 800
rect 298282 0 298338 800
rect 299294 0 299350 800
rect 300306 0 300362 800
rect 301318 0 301374 800
rect 302330 0 302386 800
rect 303342 0 303398 800
rect 304354 0 304410 800
rect 305366 0 305422 800
rect 306378 0 306434 800
rect 307390 0 307446 800
rect 308402 0 308458 800
rect 309414 0 309470 800
rect 310426 0 310482 800
rect 311438 0 311494 800
rect 312450 0 312506 800
rect 313462 0 313518 800
rect 314474 0 314530 800
rect 315486 0 315542 800
rect 316498 0 316554 800
rect 317510 0 317566 800
rect 318522 0 318578 800
rect 319534 0 319590 800
rect 320546 0 320602 800
rect 321558 0 321614 800
rect 322570 0 322626 800
rect 323582 0 323638 800
rect 324594 0 324650 800
rect 325606 0 325662 800
rect 326618 0 326674 800
rect 327630 0 327686 800
rect 328642 0 328698 800
rect 329654 0 329710 800
rect 330666 0 330722 800
rect 331678 0 331734 800
rect 332690 0 332746 800
rect 333702 0 333758 800
rect 334714 0 334770 800
rect 335726 0 335782 800
rect 336738 0 336794 800
rect 337750 0 337806 800
rect 338762 0 338818 800
rect 339774 0 339830 800
rect 340786 0 340842 800
rect 341798 0 341854 800
rect 342810 0 342866 800
rect 343822 0 343878 800
rect 344834 0 344890 800
rect 345846 0 345902 800
rect 346858 0 346914 800
rect 347870 0 347926 800
rect 348882 0 348938 800
rect 349894 0 349950 800
rect 350906 0 350962 800
rect 351918 0 351974 800
rect 352930 0 352986 800
rect 353942 0 353998 800
rect 354954 0 355010 800
rect 355966 0 356022 800
rect 356978 0 357034 800
rect 357990 0 358046 800
rect 359002 0 359058 800
rect 360014 0 360070 800
rect 361026 0 361082 800
rect 362038 0 362094 800
rect 363050 0 363106 800
rect 364062 0 364118 800
rect 365074 0 365130 800
rect 366086 0 366142 800
rect 367098 0 367154 800
rect 368110 0 368166 800
rect 369122 0 369178 800
rect 370134 0 370190 800
rect 371146 0 371202 800
rect 372158 0 372214 800
rect 373170 0 373226 800
rect 374182 0 374238 800
rect 375194 0 375250 800
rect 376206 0 376262 800
rect 377218 0 377274 800
rect 378230 0 378286 800
rect 379242 0 379298 800
rect 380254 0 380310 800
rect 381266 0 381322 800
rect 382278 0 382334 800
rect 383290 0 383346 800
rect 384302 0 384358 800
rect 385314 0 385370 800
rect 386326 0 386382 800
rect 387338 0 387394 800
rect 388350 0 388406 800
rect 389362 0 389418 800
rect 390374 0 390430 800
rect 391386 0 391442 800
rect 392398 0 392454 800
rect 393410 0 393466 800
rect 394422 0 394478 800
rect 395434 0 395490 800
rect 396446 0 396502 800
rect 397458 0 397514 800
rect 398470 0 398526 800
rect 399482 0 399538 800
rect 400494 0 400550 800
rect 401506 0 401562 800
rect 402518 0 402574 800
rect 403530 0 403586 800
rect 404542 0 404598 800
rect 405554 0 405610 800
rect 406566 0 406622 800
rect 407578 0 407634 800
rect 408590 0 408646 800
rect 409602 0 409658 800
rect 410614 0 410670 800
rect 411626 0 411682 800
rect 412638 0 412694 800
rect 413650 0 413706 800
rect 414662 0 414718 800
rect 415674 0 415730 800
rect 416686 0 416742 800
rect 417698 0 417754 800
rect 418710 0 418766 800
rect 419722 0 419778 800
rect 420734 0 420790 800
rect 421746 0 421802 800
rect 422758 0 422814 800
rect 423770 0 423826 800
rect 424782 0 424838 800
rect 425794 0 425850 800
rect 426806 0 426862 800
rect 427818 0 427874 800
rect 428830 0 428886 800
rect 429842 0 429898 800
rect 430854 0 430910 800
rect 431866 0 431922 800
rect 432878 0 432934 800
rect 433890 0 433946 800
rect 434902 0 434958 800
rect 435914 0 435970 800
rect 436926 0 436982 800
rect 437938 0 437994 800
rect 438950 0 439006 800
rect 439962 0 440018 800
rect 440974 0 441030 800
rect 441986 0 442042 800
rect 442998 0 443054 800
rect 444010 0 444066 800
rect 445022 0 445078 800
rect 446034 0 446090 800
rect 447046 0 447102 800
rect 448058 0 448114 800
rect 449070 0 449126 800
rect 450082 0 450138 800
rect 451094 0 451150 800
rect 452106 0 452162 800
rect 453118 0 453174 800
rect 454130 0 454186 800
rect 455142 0 455198 800
rect 456154 0 456210 800
rect 457166 0 457222 800
rect 458178 0 458234 800
rect 459190 0 459246 800
rect 460202 0 460258 800
rect 461214 0 461270 800
rect 462226 0 462282 800
rect 463238 0 463294 800
rect 464250 0 464306 800
rect 465262 0 465318 800
rect 466274 0 466330 800
rect 467286 0 467342 800
rect 468298 0 468354 800
rect 469310 0 469366 800
rect 470322 0 470378 800
rect 471334 0 471390 800
rect 472346 0 472402 800
rect 473358 0 473414 800
rect 474370 0 474426 800
rect 475382 0 475438 800
rect 476394 0 476450 800
rect 477406 0 477462 800
rect 478418 0 478474 800
rect 479430 0 479486 800
rect 480442 0 480498 800
rect 481454 0 481510 800
rect 482466 0 482522 800
rect 483478 0 483534 800
rect 484490 0 484546 800
rect 485502 0 485558 800
rect 486514 0 486570 800
rect 487526 0 487582 800
rect 488538 0 488594 800
rect 489550 0 489606 800
rect 490562 0 490618 800
rect 491574 0 491630 800
rect 492586 0 492642 800
rect 493598 0 493654 800
rect 494610 0 494666 800
rect 495622 0 495678 800
rect 496634 0 496690 800
rect 497646 0 497702 800
rect 498658 0 498714 800
rect 499670 0 499726 800
rect 500682 0 500738 800
rect 501694 0 501750 800
rect 502706 0 502762 800
rect 503718 0 503774 800
rect 504730 0 504786 800
rect 505742 0 505798 800
rect 506754 0 506810 800
rect 507766 0 507822 800
rect 508778 0 508834 800
rect 509790 0 509846 800
rect 510802 0 510858 800
rect 511814 0 511870 800
rect 512826 0 512882 800
rect 513838 0 513894 800
rect 514850 0 514906 800
rect 515862 0 515918 800
rect 516874 0 516930 800
rect 517886 0 517942 800
rect 518898 0 518954 800
<< obsm2 >>
rect 938 319144 10358 319200
rect 10526 319144 30322 319200
rect 30490 319144 50286 319200
rect 50454 319144 70250 319200
rect 70418 319144 90214 319200
rect 90382 319144 110178 319200
rect 110346 319144 130142 319200
rect 130310 319144 150106 319200
rect 150274 319144 170070 319200
rect 170238 319144 190034 319200
rect 190202 319144 209998 319200
rect 210166 319144 229962 319200
rect 230130 319144 249926 319200
rect 250094 319144 269890 319200
rect 270058 319144 289854 319200
rect 290022 319144 309818 319200
rect 309986 319144 329782 319200
rect 329950 319144 349746 319200
rect 349914 319144 369710 319200
rect 369878 319144 389674 319200
rect 389842 319144 409638 319200
rect 409806 319144 429602 319200
rect 429770 319144 449566 319200
rect 449734 319144 469530 319200
rect 469698 319144 489494 319200
rect 489662 319144 509458 319200
rect 509626 319144 529422 319200
rect 529590 319144 539010 319200
rect 938 856 539010 319144
rect 938 70 20938 856
rect 21106 70 21950 856
rect 22118 70 22962 856
rect 23130 70 23974 856
rect 24142 70 24986 856
rect 25154 70 25998 856
rect 26166 70 27010 856
rect 27178 70 28022 856
rect 28190 70 29034 856
rect 29202 70 30046 856
rect 30214 70 31058 856
rect 31226 70 32070 856
rect 32238 70 33082 856
rect 33250 70 34094 856
rect 34262 70 35106 856
rect 35274 70 36118 856
rect 36286 70 37130 856
rect 37298 70 38142 856
rect 38310 70 39154 856
rect 39322 70 40166 856
rect 40334 70 41178 856
rect 41346 70 42190 856
rect 42358 70 43202 856
rect 43370 70 44214 856
rect 44382 70 45226 856
rect 45394 70 46238 856
rect 46406 70 47250 856
rect 47418 70 48262 856
rect 48430 70 49274 856
rect 49442 70 50286 856
rect 50454 70 51298 856
rect 51466 70 52310 856
rect 52478 70 53322 856
rect 53490 70 54334 856
rect 54502 70 55346 856
rect 55514 70 56358 856
rect 56526 70 57370 856
rect 57538 70 58382 856
rect 58550 70 59394 856
rect 59562 70 60406 856
rect 60574 70 61418 856
rect 61586 70 62430 856
rect 62598 70 63442 856
rect 63610 70 64454 856
rect 64622 70 65466 856
rect 65634 70 66478 856
rect 66646 70 67490 856
rect 67658 70 68502 856
rect 68670 70 69514 856
rect 69682 70 70526 856
rect 70694 70 71538 856
rect 71706 70 72550 856
rect 72718 70 73562 856
rect 73730 70 74574 856
rect 74742 70 75586 856
rect 75754 70 76598 856
rect 76766 70 77610 856
rect 77778 70 78622 856
rect 78790 70 79634 856
rect 79802 70 80646 856
rect 80814 70 81658 856
rect 81826 70 82670 856
rect 82838 70 83682 856
rect 83850 70 84694 856
rect 84862 70 85706 856
rect 85874 70 86718 856
rect 86886 70 87730 856
rect 87898 70 88742 856
rect 88910 70 89754 856
rect 89922 70 90766 856
rect 90934 70 91778 856
rect 91946 70 92790 856
rect 92958 70 93802 856
rect 93970 70 94814 856
rect 94982 70 95826 856
rect 95994 70 96838 856
rect 97006 70 97850 856
rect 98018 70 98862 856
rect 99030 70 99874 856
rect 100042 70 100886 856
rect 101054 70 101898 856
rect 102066 70 102910 856
rect 103078 70 103922 856
rect 104090 70 104934 856
rect 105102 70 105946 856
rect 106114 70 106958 856
rect 107126 70 107970 856
rect 108138 70 108982 856
rect 109150 70 109994 856
rect 110162 70 111006 856
rect 111174 70 112018 856
rect 112186 70 113030 856
rect 113198 70 114042 856
rect 114210 70 115054 856
rect 115222 70 116066 856
rect 116234 70 117078 856
rect 117246 70 118090 856
rect 118258 70 119102 856
rect 119270 70 120114 856
rect 120282 70 121126 856
rect 121294 70 122138 856
rect 122306 70 123150 856
rect 123318 70 124162 856
rect 124330 70 125174 856
rect 125342 70 126186 856
rect 126354 70 127198 856
rect 127366 70 128210 856
rect 128378 70 129222 856
rect 129390 70 130234 856
rect 130402 70 131246 856
rect 131414 70 132258 856
rect 132426 70 133270 856
rect 133438 70 134282 856
rect 134450 70 135294 856
rect 135462 70 136306 856
rect 136474 70 137318 856
rect 137486 70 138330 856
rect 138498 70 139342 856
rect 139510 70 140354 856
rect 140522 70 141366 856
rect 141534 70 142378 856
rect 142546 70 143390 856
rect 143558 70 144402 856
rect 144570 70 145414 856
rect 145582 70 146426 856
rect 146594 70 147438 856
rect 147606 70 148450 856
rect 148618 70 149462 856
rect 149630 70 150474 856
rect 150642 70 151486 856
rect 151654 70 152498 856
rect 152666 70 153510 856
rect 153678 70 154522 856
rect 154690 70 155534 856
rect 155702 70 156546 856
rect 156714 70 157558 856
rect 157726 70 158570 856
rect 158738 70 159582 856
rect 159750 70 160594 856
rect 160762 70 161606 856
rect 161774 70 162618 856
rect 162786 70 163630 856
rect 163798 70 164642 856
rect 164810 70 165654 856
rect 165822 70 166666 856
rect 166834 70 167678 856
rect 167846 70 168690 856
rect 168858 70 169702 856
rect 169870 70 170714 856
rect 170882 70 171726 856
rect 171894 70 172738 856
rect 172906 70 173750 856
rect 173918 70 174762 856
rect 174930 70 175774 856
rect 175942 70 176786 856
rect 176954 70 177798 856
rect 177966 70 178810 856
rect 178978 70 179822 856
rect 179990 70 180834 856
rect 181002 70 181846 856
rect 182014 70 182858 856
rect 183026 70 183870 856
rect 184038 70 184882 856
rect 185050 70 185894 856
rect 186062 70 186906 856
rect 187074 70 187918 856
rect 188086 70 188930 856
rect 189098 70 189942 856
rect 190110 70 190954 856
rect 191122 70 191966 856
rect 192134 70 192978 856
rect 193146 70 193990 856
rect 194158 70 195002 856
rect 195170 70 196014 856
rect 196182 70 197026 856
rect 197194 70 198038 856
rect 198206 70 199050 856
rect 199218 70 200062 856
rect 200230 70 201074 856
rect 201242 70 202086 856
rect 202254 70 203098 856
rect 203266 70 204110 856
rect 204278 70 205122 856
rect 205290 70 206134 856
rect 206302 70 207146 856
rect 207314 70 208158 856
rect 208326 70 209170 856
rect 209338 70 210182 856
rect 210350 70 211194 856
rect 211362 70 212206 856
rect 212374 70 213218 856
rect 213386 70 214230 856
rect 214398 70 215242 856
rect 215410 70 216254 856
rect 216422 70 217266 856
rect 217434 70 218278 856
rect 218446 70 219290 856
rect 219458 70 220302 856
rect 220470 70 221314 856
rect 221482 70 222326 856
rect 222494 70 223338 856
rect 223506 70 224350 856
rect 224518 70 225362 856
rect 225530 70 226374 856
rect 226542 70 227386 856
rect 227554 70 228398 856
rect 228566 70 229410 856
rect 229578 70 230422 856
rect 230590 70 231434 856
rect 231602 70 232446 856
rect 232614 70 233458 856
rect 233626 70 234470 856
rect 234638 70 235482 856
rect 235650 70 236494 856
rect 236662 70 237506 856
rect 237674 70 238518 856
rect 238686 70 239530 856
rect 239698 70 240542 856
rect 240710 70 241554 856
rect 241722 70 242566 856
rect 242734 70 243578 856
rect 243746 70 244590 856
rect 244758 70 245602 856
rect 245770 70 246614 856
rect 246782 70 247626 856
rect 247794 70 248638 856
rect 248806 70 249650 856
rect 249818 70 250662 856
rect 250830 70 251674 856
rect 251842 70 252686 856
rect 252854 70 253698 856
rect 253866 70 254710 856
rect 254878 70 255722 856
rect 255890 70 256734 856
rect 256902 70 257746 856
rect 257914 70 258758 856
rect 258926 70 259770 856
rect 259938 70 260782 856
rect 260950 70 261794 856
rect 261962 70 262806 856
rect 262974 70 263818 856
rect 263986 70 264830 856
rect 264998 70 265842 856
rect 266010 70 266854 856
rect 267022 70 267866 856
rect 268034 70 268878 856
rect 269046 70 269890 856
rect 270058 70 270902 856
rect 271070 70 271914 856
rect 272082 70 272926 856
rect 273094 70 273938 856
rect 274106 70 274950 856
rect 275118 70 275962 856
rect 276130 70 276974 856
rect 277142 70 277986 856
rect 278154 70 278998 856
rect 279166 70 280010 856
rect 280178 70 281022 856
rect 281190 70 282034 856
rect 282202 70 283046 856
rect 283214 70 284058 856
rect 284226 70 285070 856
rect 285238 70 286082 856
rect 286250 70 287094 856
rect 287262 70 288106 856
rect 288274 70 289118 856
rect 289286 70 290130 856
rect 290298 70 291142 856
rect 291310 70 292154 856
rect 292322 70 293166 856
rect 293334 70 294178 856
rect 294346 70 295190 856
rect 295358 70 296202 856
rect 296370 70 297214 856
rect 297382 70 298226 856
rect 298394 70 299238 856
rect 299406 70 300250 856
rect 300418 70 301262 856
rect 301430 70 302274 856
rect 302442 70 303286 856
rect 303454 70 304298 856
rect 304466 70 305310 856
rect 305478 70 306322 856
rect 306490 70 307334 856
rect 307502 70 308346 856
rect 308514 70 309358 856
rect 309526 70 310370 856
rect 310538 70 311382 856
rect 311550 70 312394 856
rect 312562 70 313406 856
rect 313574 70 314418 856
rect 314586 70 315430 856
rect 315598 70 316442 856
rect 316610 70 317454 856
rect 317622 70 318466 856
rect 318634 70 319478 856
rect 319646 70 320490 856
rect 320658 70 321502 856
rect 321670 70 322514 856
rect 322682 70 323526 856
rect 323694 70 324538 856
rect 324706 70 325550 856
rect 325718 70 326562 856
rect 326730 70 327574 856
rect 327742 70 328586 856
rect 328754 70 329598 856
rect 329766 70 330610 856
rect 330778 70 331622 856
rect 331790 70 332634 856
rect 332802 70 333646 856
rect 333814 70 334658 856
rect 334826 70 335670 856
rect 335838 70 336682 856
rect 336850 70 337694 856
rect 337862 70 338706 856
rect 338874 70 339718 856
rect 339886 70 340730 856
rect 340898 70 341742 856
rect 341910 70 342754 856
rect 342922 70 343766 856
rect 343934 70 344778 856
rect 344946 70 345790 856
rect 345958 70 346802 856
rect 346970 70 347814 856
rect 347982 70 348826 856
rect 348994 70 349838 856
rect 350006 70 350850 856
rect 351018 70 351862 856
rect 352030 70 352874 856
rect 353042 70 353886 856
rect 354054 70 354898 856
rect 355066 70 355910 856
rect 356078 70 356922 856
rect 357090 70 357934 856
rect 358102 70 358946 856
rect 359114 70 359958 856
rect 360126 70 360970 856
rect 361138 70 361982 856
rect 362150 70 362994 856
rect 363162 70 364006 856
rect 364174 70 365018 856
rect 365186 70 366030 856
rect 366198 70 367042 856
rect 367210 70 368054 856
rect 368222 70 369066 856
rect 369234 70 370078 856
rect 370246 70 371090 856
rect 371258 70 372102 856
rect 372270 70 373114 856
rect 373282 70 374126 856
rect 374294 70 375138 856
rect 375306 70 376150 856
rect 376318 70 377162 856
rect 377330 70 378174 856
rect 378342 70 379186 856
rect 379354 70 380198 856
rect 380366 70 381210 856
rect 381378 70 382222 856
rect 382390 70 383234 856
rect 383402 70 384246 856
rect 384414 70 385258 856
rect 385426 70 386270 856
rect 386438 70 387282 856
rect 387450 70 388294 856
rect 388462 70 389306 856
rect 389474 70 390318 856
rect 390486 70 391330 856
rect 391498 70 392342 856
rect 392510 70 393354 856
rect 393522 70 394366 856
rect 394534 70 395378 856
rect 395546 70 396390 856
rect 396558 70 397402 856
rect 397570 70 398414 856
rect 398582 70 399426 856
rect 399594 70 400438 856
rect 400606 70 401450 856
rect 401618 70 402462 856
rect 402630 70 403474 856
rect 403642 70 404486 856
rect 404654 70 405498 856
rect 405666 70 406510 856
rect 406678 70 407522 856
rect 407690 70 408534 856
rect 408702 70 409546 856
rect 409714 70 410558 856
rect 410726 70 411570 856
rect 411738 70 412582 856
rect 412750 70 413594 856
rect 413762 70 414606 856
rect 414774 70 415618 856
rect 415786 70 416630 856
rect 416798 70 417642 856
rect 417810 70 418654 856
rect 418822 70 419666 856
rect 419834 70 420678 856
rect 420846 70 421690 856
rect 421858 70 422702 856
rect 422870 70 423714 856
rect 423882 70 424726 856
rect 424894 70 425738 856
rect 425906 70 426750 856
rect 426918 70 427762 856
rect 427930 70 428774 856
rect 428942 70 429786 856
rect 429954 70 430798 856
rect 430966 70 431810 856
rect 431978 70 432822 856
rect 432990 70 433834 856
rect 434002 70 434846 856
rect 435014 70 435858 856
rect 436026 70 436870 856
rect 437038 70 437882 856
rect 438050 70 438894 856
rect 439062 70 439906 856
rect 440074 70 440918 856
rect 441086 70 441930 856
rect 442098 70 442942 856
rect 443110 70 443954 856
rect 444122 70 444966 856
rect 445134 70 445978 856
rect 446146 70 446990 856
rect 447158 70 448002 856
rect 448170 70 449014 856
rect 449182 70 450026 856
rect 450194 70 451038 856
rect 451206 70 452050 856
rect 452218 70 453062 856
rect 453230 70 454074 856
rect 454242 70 455086 856
rect 455254 70 456098 856
rect 456266 70 457110 856
rect 457278 70 458122 856
rect 458290 70 459134 856
rect 459302 70 460146 856
rect 460314 70 461158 856
rect 461326 70 462170 856
rect 462338 70 463182 856
rect 463350 70 464194 856
rect 464362 70 465206 856
rect 465374 70 466218 856
rect 466386 70 467230 856
rect 467398 70 468242 856
rect 468410 70 469254 856
rect 469422 70 470266 856
rect 470434 70 471278 856
rect 471446 70 472290 856
rect 472458 70 473302 856
rect 473470 70 474314 856
rect 474482 70 475326 856
rect 475494 70 476338 856
rect 476506 70 477350 856
rect 477518 70 478362 856
rect 478530 70 479374 856
rect 479542 70 480386 856
rect 480554 70 481398 856
rect 481566 70 482410 856
rect 482578 70 483422 856
rect 483590 70 484434 856
rect 484602 70 485446 856
rect 485614 70 486458 856
rect 486626 70 487470 856
rect 487638 70 488482 856
rect 488650 70 489494 856
rect 489662 70 490506 856
rect 490674 70 491518 856
rect 491686 70 492530 856
rect 492698 70 493542 856
rect 493710 70 494554 856
rect 494722 70 495566 856
rect 495734 70 496578 856
rect 496746 70 497590 856
rect 497758 70 498602 856
rect 498770 70 499614 856
rect 499782 70 500626 856
rect 500794 70 501638 856
rect 501806 70 502650 856
rect 502818 70 503662 856
rect 503830 70 504674 856
rect 504842 70 505686 856
rect 505854 70 506698 856
rect 506866 70 507710 856
rect 507878 70 508722 856
rect 508890 70 509734 856
rect 509902 70 510746 856
rect 510914 70 511758 856
rect 511926 70 512770 856
rect 512938 70 513782 856
rect 513950 70 514794 856
rect 514962 70 515806 856
rect 515974 70 516818 856
rect 516986 70 517830 856
rect 517998 70 518842 856
rect 519010 70 539010 856
<< metal3 >>
rect 0 316072 800 316192
rect 539200 315528 540000 315648
rect 0 308456 800 308576
rect 539200 308456 540000 308576
rect 539200 301384 540000 301504
rect 0 300840 800 300960
rect 539200 294312 540000 294432
rect 0 293224 800 293344
rect 539200 287240 540000 287360
rect 0 285608 800 285728
rect 539200 280168 540000 280288
rect 0 277992 800 278112
rect 539200 273096 540000 273216
rect 0 270376 800 270496
rect 539200 266024 540000 266144
rect 0 262760 800 262880
rect 539200 258952 540000 259072
rect 0 255144 800 255264
rect 539200 251880 540000 252000
rect 0 247528 800 247648
rect 539200 244808 540000 244928
rect 0 239912 800 240032
rect 539200 237736 540000 237856
rect 0 232296 800 232416
rect 539200 230664 540000 230784
rect 0 224680 800 224800
rect 539200 223592 540000 223712
rect 0 217064 800 217184
rect 539200 216520 540000 216640
rect 0 209448 800 209568
rect 539200 209448 540000 209568
rect 539200 202376 540000 202496
rect 0 201832 800 201952
rect 539200 195304 540000 195424
rect 0 194216 800 194336
rect 539200 188232 540000 188352
rect 0 186600 800 186720
rect 539200 181160 540000 181280
rect 0 178984 800 179104
rect 539200 174088 540000 174208
rect 0 171368 800 171488
rect 539200 167016 540000 167136
rect 0 163752 800 163872
rect 539200 159944 540000 160064
rect 0 156136 800 156256
rect 539200 152872 540000 152992
rect 0 148520 800 148640
rect 539200 145800 540000 145920
rect 0 140904 800 141024
rect 539200 138728 540000 138848
rect 0 133288 800 133408
rect 539200 131656 540000 131776
rect 0 125672 800 125792
rect 539200 124584 540000 124704
rect 0 118056 800 118176
rect 539200 117512 540000 117632
rect 0 110440 800 110560
rect 539200 110440 540000 110560
rect 539200 103368 540000 103488
rect 0 102824 800 102944
rect 539200 96296 540000 96416
rect 0 95208 800 95328
rect 539200 89224 540000 89344
rect 0 87592 800 87712
rect 539200 82152 540000 82272
rect 0 79976 800 80096
rect 539200 75080 540000 75200
rect 0 72360 800 72480
rect 539200 68008 540000 68128
rect 0 64744 800 64864
rect 539200 60936 540000 61056
rect 0 57128 800 57248
rect 539200 53864 540000 53984
rect 0 49512 800 49632
rect 539200 46792 540000 46912
rect 0 41896 800 42016
rect 539200 39720 540000 39840
rect 0 34280 800 34400
rect 539200 32648 540000 32768
rect 0 26664 800 26784
rect 539200 25576 540000 25696
rect 0 19048 800 19168
rect 539200 18504 540000 18624
rect 0 11432 800 11552
rect 539200 11432 540000 11552
rect 539200 4360 540000 4480
rect 0 3816 800 3936
<< obsm3 >>
rect 798 316272 539200 317729
rect 880 315992 539200 316272
rect 798 315728 539200 315992
rect 798 315448 539120 315728
rect 798 308656 539200 315448
rect 880 308376 539120 308656
rect 798 301584 539200 308376
rect 798 301304 539120 301584
rect 798 301040 539200 301304
rect 880 300760 539200 301040
rect 798 294512 539200 300760
rect 798 294232 539120 294512
rect 798 293424 539200 294232
rect 880 293144 539200 293424
rect 798 287440 539200 293144
rect 798 287160 539120 287440
rect 798 285808 539200 287160
rect 880 285528 539200 285808
rect 798 280368 539200 285528
rect 798 280088 539120 280368
rect 798 278192 539200 280088
rect 880 277912 539200 278192
rect 798 273296 539200 277912
rect 798 273016 539120 273296
rect 798 270576 539200 273016
rect 880 270296 539200 270576
rect 798 266224 539200 270296
rect 798 265944 539120 266224
rect 798 262960 539200 265944
rect 880 262680 539200 262960
rect 798 259152 539200 262680
rect 798 258872 539120 259152
rect 798 255344 539200 258872
rect 880 255064 539200 255344
rect 798 252080 539200 255064
rect 798 251800 539120 252080
rect 798 247728 539200 251800
rect 880 247448 539200 247728
rect 798 245008 539200 247448
rect 798 244728 539120 245008
rect 798 240112 539200 244728
rect 880 239832 539200 240112
rect 798 237936 539200 239832
rect 798 237656 539120 237936
rect 798 232496 539200 237656
rect 880 232216 539200 232496
rect 798 230864 539200 232216
rect 798 230584 539120 230864
rect 798 224880 539200 230584
rect 880 224600 539200 224880
rect 798 223792 539200 224600
rect 798 223512 539120 223792
rect 798 217264 539200 223512
rect 880 216984 539200 217264
rect 798 216720 539200 216984
rect 798 216440 539120 216720
rect 798 209648 539200 216440
rect 880 209368 539120 209648
rect 798 202576 539200 209368
rect 798 202296 539120 202576
rect 798 202032 539200 202296
rect 880 201752 539200 202032
rect 798 195504 539200 201752
rect 798 195224 539120 195504
rect 798 194416 539200 195224
rect 880 194136 539200 194416
rect 798 188432 539200 194136
rect 798 188152 539120 188432
rect 798 186800 539200 188152
rect 880 186520 539200 186800
rect 798 181360 539200 186520
rect 798 181080 539120 181360
rect 798 179184 539200 181080
rect 880 178904 539200 179184
rect 798 174288 539200 178904
rect 798 174008 539120 174288
rect 798 171568 539200 174008
rect 880 171288 539200 171568
rect 798 167216 539200 171288
rect 798 166936 539120 167216
rect 798 163952 539200 166936
rect 880 163672 539200 163952
rect 798 160144 539200 163672
rect 798 159864 539120 160144
rect 798 156336 539200 159864
rect 880 156056 539200 156336
rect 798 153072 539200 156056
rect 798 152792 539120 153072
rect 798 148720 539200 152792
rect 880 148440 539200 148720
rect 798 146000 539200 148440
rect 798 145720 539120 146000
rect 798 141104 539200 145720
rect 880 140824 539200 141104
rect 798 138928 539200 140824
rect 798 138648 539120 138928
rect 798 133488 539200 138648
rect 880 133208 539200 133488
rect 798 131856 539200 133208
rect 798 131576 539120 131856
rect 798 125872 539200 131576
rect 880 125592 539200 125872
rect 798 124784 539200 125592
rect 798 124504 539120 124784
rect 798 118256 539200 124504
rect 880 117976 539200 118256
rect 798 117712 539200 117976
rect 798 117432 539120 117712
rect 798 110640 539200 117432
rect 880 110360 539120 110640
rect 798 103568 539200 110360
rect 798 103288 539120 103568
rect 798 103024 539200 103288
rect 880 102744 539200 103024
rect 798 96496 539200 102744
rect 798 96216 539120 96496
rect 798 95408 539200 96216
rect 880 95128 539200 95408
rect 798 89424 539200 95128
rect 798 89144 539120 89424
rect 798 87792 539200 89144
rect 880 87512 539200 87792
rect 798 82352 539200 87512
rect 798 82072 539120 82352
rect 798 80176 539200 82072
rect 880 79896 539200 80176
rect 798 75280 539200 79896
rect 798 75000 539120 75280
rect 798 72560 539200 75000
rect 880 72280 539200 72560
rect 798 68208 539200 72280
rect 798 67928 539120 68208
rect 798 64944 539200 67928
rect 880 64664 539200 64944
rect 798 61136 539200 64664
rect 798 60856 539120 61136
rect 798 57328 539200 60856
rect 880 57048 539200 57328
rect 798 54064 539200 57048
rect 798 53784 539120 54064
rect 798 49712 539200 53784
rect 880 49432 539200 49712
rect 798 46992 539200 49432
rect 798 46712 539120 46992
rect 798 42096 539200 46712
rect 880 41816 539200 42096
rect 798 39920 539200 41816
rect 798 39640 539120 39920
rect 798 34480 539200 39640
rect 880 34200 539200 34480
rect 798 32848 539200 34200
rect 798 32568 539120 32848
rect 798 26864 539200 32568
rect 880 26584 539200 26864
rect 798 25776 539200 26584
rect 798 25496 539120 25776
rect 798 19248 539200 25496
rect 880 18968 539200 19248
rect 798 18704 539200 18968
rect 798 18424 539120 18704
rect 798 11632 539200 18424
rect 880 11352 539120 11632
rect 798 4560 539200 11352
rect 798 4280 539120 4560
rect 798 4016 539200 4280
rect 880 3736 539200 4016
rect 798 1803 539200 3736
<< metal4 >>
rect 4208 2128 4528 317744
rect 19568 2128 19888 317744
rect 34928 2128 35248 317744
rect 50288 2128 50608 317744
rect 65648 2128 65968 317744
rect 81008 2128 81328 317744
rect 96368 2128 96688 317744
rect 111728 2128 112048 317744
rect 127088 2128 127408 317744
rect 142448 2128 142768 317744
rect 157808 2128 158128 317744
rect 173168 2128 173488 317744
rect 188528 2128 188848 317744
rect 203888 2128 204208 317744
rect 219248 2128 219568 317744
rect 234608 2128 234928 317744
rect 249968 2128 250288 317744
rect 265328 2128 265648 317744
rect 280688 2128 281008 317744
rect 296048 2128 296368 317744
rect 311408 2128 311728 317744
rect 326768 2128 327088 317744
rect 342128 2128 342448 317744
rect 357488 2128 357808 317744
rect 372848 2128 373168 317744
rect 388208 2128 388528 317744
rect 403568 2128 403888 317744
rect 418928 2128 419248 317744
rect 434288 2128 434608 317744
rect 449648 2128 449968 317744
rect 465008 2128 465328 317744
rect 480368 2128 480688 317744
rect 495728 2128 496048 317744
rect 511088 2128 511408 317744
rect 526448 2128 526768 317744
<< obsm4 >>
rect 235027 3299 249888 84149
rect 250368 3299 265248 84149
rect 265728 3299 280608 84149
rect 281088 3299 295968 84149
rect 296448 3299 311328 84149
rect 311808 3299 326688 84149
rect 327168 3299 342048 84149
rect 342528 3299 357408 84149
rect 357888 3299 367389 84149
<< labels >>
rlabel metal3 s 539200 4360 540000 4480 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 539200 216520 540000 216640 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 539200 237736 540000 237856 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 539200 258952 540000 259072 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 539200 280168 540000 280288 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 539200 301384 540000 301504 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 529478 319200 529534 320000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 469586 319200 469642 320000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 409694 319200 409750 320000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 349802 319200 349858 320000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 289910 319200 289966 320000 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 539200 25576 540000 25696 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 230018 319200 230074 320000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 170126 319200 170182 320000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 110234 319200 110290 320000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 50342 319200 50398 320000 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s 0 316072 800 316192 6 io_in[24]
port 17 nsew signal input
rlabel metal3 s 0 293224 800 293344 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 0 270376 800 270496 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 0 247528 800 247648 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 0 224680 800 224800 6 io_in[28]
port 21 nsew signal input
rlabel metal3 s 0 201832 800 201952 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 539200 46792 540000 46912 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s 0 178984 800 179104 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 0 156136 800 156256 6 io_in[31]
port 25 nsew signal input
rlabel metal3 s 0 133288 800 133408 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 0 110440 800 110560 6 io_in[33]
port 27 nsew signal input
rlabel metal3 s 0 87592 800 87712 6 io_in[34]
port 28 nsew signal input
rlabel metal3 s 0 64744 800 64864 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 0 41896 800 42016 6 io_in[36]
port 30 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 539200 68008 540000 68128 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 539200 89224 540000 89344 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 539200 110440 540000 110560 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 539200 131656 540000 131776 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 539200 152872 540000 152992 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 539200 174088 540000 174208 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 539200 195304 540000 195424 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 539200 18504 540000 18624 6 io_oeb[0]
port 39 nsew signal output
rlabel metal3 s 539200 230664 540000 230784 6 io_oeb[10]
port 40 nsew signal output
rlabel metal3 s 539200 251880 540000 252000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal3 s 539200 273096 540000 273216 6 io_oeb[12]
port 42 nsew signal output
rlabel metal3 s 539200 294312 540000 294432 6 io_oeb[13]
port 43 nsew signal output
rlabel metal3 s 539200 315528 540000 315648 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 489550 319200 489606 320000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 429658 319200 429714 320000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 369766 319200 369822 320000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 309874 319200 309930 320000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 249982 319200 250038 320000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal3 s 539200 39720 540000 39840 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 190090 319200 190146 320000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 130198 319200 130254 320000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 70306 319200 70362 320000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 10414 319200 10470 320000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s 0 300840 800 300960 6 io_oeb[24]
port 55 nsew signal output
rlabel metal3 s 0 277992 800 278112 6 io_oeb[25]
port 56 nsew signal output
rlabel metal3 s 0 255144 800 255264 6 io_oeb[26]
port 57 nsew signal output
rlabel metal3 s 0 232296 800 232416 6 io_oeb[27]
port 58 nsew signal output
rlabel metal3 s 0 209448 800 209568 6 io_oeb[28]
port 59 nsew signal output
rlabel metal3 s 0 186600 800 186720 6 io_oeb[29]
port 60 nsew signal output
rlabel metal3 s 539200 60936 540000 61056 6 io_oeb[2]
port 61 nsew signal output
rlabel metal3 s 0 163752 800 163872 6 io_oeb[30]
port 62 nsew signal output
rlabel metal3 s 0 140904 800 141024 6 io_oeb[31]
port 63 nsew signal output
rlabel metal3 s 0 118056 800 118176 6 io_oeb[32]
port 64 nsew signal output
rlabel metal3 s 0 95208 800 95328 6 io_oeb[33]
port 65 nsew signal output
rlabel metal3 s 0 72360 800 72480 6 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s 0 49512 800 49632 6 io_oeb[35]
port 67 nsew signal output
rlabel metal3 s 0 26664 800 26784 6 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s 0 3816 800 3936 6 io_oeb[37]
port 69 nsew signal output
rlabel metal3 s 539200 82152 540000 82272 6 io_oeb[3]
port 70 nsew signal output
rlabel metal3 s 539200 103368 540000 103488 6 io_oeb[4]
port 71 nsew signal output
rlabel metal3 s 539200 124584 540000 124704 6 io_oeb[5]
port 72 nsew signal output
rlabel metal3 s 539200 145800 540000 145920 6 io_oeb[6]
port 73 nsew signal output
rlabel metal3 s 539200 167016 540000 167136 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 539200 188232 540000 188352 6 io_oeb[8]
port 75 nsew signal output
rlabel metal3 s 539200 209448 540000 209568 6 io_oeb[9]
port 76 nsew signal output
rlabel metal3 s 539200 11432 540000 11552 6 io_out[0]
port 77 nsew signal output
rlabel metal3 s 539200 223592 540000 223712 6 io_out[10]
port 78 nsew signal output
rlabel metal3 s 539200 244808 540000 244928 6 io_out[11]
port 79 nsew signal output
rlabel metal3 s 539200 266024 540000 266144 6 io_out[12]
port 80 nsew signal output
rlabel metal3 s 539200 287240 540000 287360 6 io_out[13]
port 81 nsew signal output
rlabel metal3 s 539200 308456 540000 308576 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 509514 319200 509570 320000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 449622 319200 449678 320000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 389730 319200 389786 320000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 329838 319200 329894 320000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 269946 319200 270002 320000 6 io_out[19]
port 87 nsew signal output
rlabel metal3 s 539200 32648 540000 32768 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 210054 319200 210110 320000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 150162 319200 150218 320000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 90270 319200 90326 320000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 30378 319200 30434 320000 6 io_out[23]
port 92 nsew signal output
rlabel metal3 s 0 308456 800 308576 6 io_out[24]
port 93 nsew signal output
rlabel metal3 s 0 285608 800 285728 6 io_out[25]
port 94 nsew signal output
rlabel metal3 s 0 262760 800 262880 6 io_out[26]
port 95 nsew signal output
rlabel metal3 s 0 239912 800 240032 6 io_out[27]
port 96 nsew signal output
rlabel metal3 s 0 217064 800 217184 6 io_out[28]
port 97 nsew signal output
rlabel metal3 s 0 194216 800 194336 6 io_out[29]
port 98 nsew signal output
rlabel metal3 s 539200 53864 540000 53984 6 io_out[2]
port 99 nsew signal output
rlabel metal3 s 0 171368 800 171488 6 io_out[30]
port 100 nsew signal output
rlabel metal3 s 0 148520 800 148640 6 io_out[31]
port 101 nsew signal output
rlabel metal3 s 0 125672 800 125792 6 io_out[32]
port 102 nsew signal output
rlabel metal3 s 0 102824 800 102944 6 io_out[33]
port 103 nsew signal output
rlabel metal3 s 0 79976 800 80096 6 io_out[34]
port 104 nsew signal output
rlabel metal3 s 0 57128 800 57248 6 io_out[35]
port 105 nsew signal output
rlabel metal3 s 0 34280 800 34400 6 io_out[36]
port 106 nsew signal output
rlabel metal3 s 0 11432 800 11552 6 io_out[37]
port 107 nsew signal output
rlabel metal3 s 539200 75080 540000 75200 6 io_out[3]
port 108 nsew signal output
rlabel metal3 s 539200 96296 540000 96416 6 io_out[4]
port 109 nsew signal output
rlabel metal3 s 539200 117512 540000 117632 6 io_out[5]
port 110 nsew signal output
rlabel metal3 s 539200 138728 540000 138848 6 io_out[6]
port 111 nsew signal output
rlabel metal3 s 539200 159944 540000 160064 6 io_out[7]
port 112 nsew signal output
rlabel metal3 s 539200 181160 540000 181280 6 io_out[8]
port 113 nsew signal output
rlabel metal3 s 539200 202376 540000 202496 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 516874 0 516930 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 517886 0 517942 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 518898 0 518954 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 128266 0 128322 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 431866 0 431922 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 434902 0 434958 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 437938 0 437994 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 440974 0 441030 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 444010 0 444066 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 447046 0 447102 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 450082 0 450138 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 453118 0 453174 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 456154 0 456210 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 459190 0 459246 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 158626 0 158682 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 462226 0 462282 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 465262 0 465318 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 468298 0 468354 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 471334 0 471390 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 474370 0 474426 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 477406 0 477462 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 480442 0 480498 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 483478 0 483534 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 486514 0 486570 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 489550 0 489606 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 161662 0 161718 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 492586 0 492642 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 495622 0 495678 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 498658 0 498714 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 501694 0 501750 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 504730 0 504786 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 507766 0 507822 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 510802 0 510858 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 513838 0 513894 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 164698 0 164754 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 167734 0 167790 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 170770 0 170826 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 173806 0 173862 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 176842 0 176898 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 179878 0 179934 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 182914 0 182970 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 185950 0 186006 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 131302 0 131358 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 188986 0 189042 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 192022 0 192078 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 195058 0 195114 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 198094 0 198150 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 201130 0 201186 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 204166 0 204222 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 207202 0 207258 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 210238 0 210294 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 213274 0 213330 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 216310 0 216366 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 134338 0 134394 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 219346 0 219402 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 222382 0 222438 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 225418 0 225474 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 228454 0 228510 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 231490 0 231546 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 234526 0 234582 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 237562 0 237618 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 240598 0 240654 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 243634 0 243690 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 246670 0 246726 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 137374 0 137430 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 249706 0 249762 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 252742 0 252798 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 255778 0 255834 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 258814 0 258870 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 261850 0 261906 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 264886 0 264942 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 267922 0 267978 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 270958 0 271014 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 273994 0 274050 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 277030 0 277086 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 140410 0 140466 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 280066 0 280122 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 283102 0 283158 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 286138 0 286194 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 289174 0 289230 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 292210 0 292266 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 295246 0 295302 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 298282 0 298338 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 301318 0 301374 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 304354 0 304410 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 307390 0 307446 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 143446 0 143502 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 310426 0 310482 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 313462 0 313518 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 316498 0 316554 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 319534 0 319590 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 322570 0 322626 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 325606 0 325662 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 328642 0 328698 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 331678 0 331734 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 334714 0 334770 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 337750 0 337806 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 146482 0 146538 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 340786 0 340842 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 343822 0 343878 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 346858 0 346914 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 349894 0 349950 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 352930 0 352986 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 355966 0 356022 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 359002 0 359058 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 362038 0 362094 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 365074 0 365130 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 368110 0 368166 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 149518 0 149574 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 371146 0 371202 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 374182 0 374238 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 377218 0 377274 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 380254 0 380310 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 383290 0 383346 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 386326 0 386382 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 389362 0 389418 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 392398 0 392454 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 395434 0 395490 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 398470 0 398526 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 152554 0 152610 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 401506 0 401562 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 404542 0 404598 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 407578 0 407634 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 410614 0 410670 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 413650 0 413706 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 416686 0 416742 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 419722 0 419778 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 422758 0 422814 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 425794 0 425850 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 428830 0 428886 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 155590 0 155646 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 129278 0 129334 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 432878 0 432934 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 435914 0 435970 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 438950 0 439006 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 441986 0 442042 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 445022 0 445078 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 448058 0 448114 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 451094 0 451150 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 454130 0 454186 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 457166 0 457222 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 460202 0 460258 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 159638 0 159694 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 463238 0 463294 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 466274 0 466330 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 469310 0 469366 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 472346 0 472402 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 475382 0 475438 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 478418 0 478474 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 481454 0 481510 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 484490 0 484546 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 487526 0 487582 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 490562 0 490618 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 162674 0 162730 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 493598 0 493654 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 496634 0 496690 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 499670 0 499726 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 502706 0 502762 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 505742 0 505798 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 508778 0 508834 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 511814 0 511870 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 514850 0 514906 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 165710 0 165766 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 168746 0 168802 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 171782 0 171838 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 174818 0 174874 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 177854 0 177910 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 180890 0 180946 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 183926 0 183982 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 186962 0 187018 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 132314 0 132370 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 189998 0 190054 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 193034 0 193090 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 196070 0 196126 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 199106 0 199162 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 202142 0 202198 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 205178 0 205234 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 208214 0 208270 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 211250 0 211306 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 214286 0 214342 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 217322 0 217378 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 135350 0 135406 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 220358 0 220414 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 223394 0 223450 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 226430 0 226486 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 229466 0 229522 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 232502 0 232558 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 235538 0 235594 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 238574 0 238630 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 241610 0 241666 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 244646 0 244702 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 247682 0 247738 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 138386 0 138442 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 250718 0 250774 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 253754 0 253810 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 256790 0 256846 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 259826 0 259882 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 262862 0 262918 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 265898 0 265954 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 268934 0 268990 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 271970 0 272026 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 275006 0 275062 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 278042 0 278098 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 141422 0 141478 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 281078 0 281134 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 284114 0 284170 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 287150 0 287206 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 290186 0 290242 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 293222 0 293278 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 296258 0 296314 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 299294 0 299350 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 302330 0 302386 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 305366 0 305422 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 308402 0 308458 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 144458 0 144514 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 311438 0 311494 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 314474 0 314530 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 317510 0 317566 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 320546 0 320602 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 323582 0 323638 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 326618 0 326674 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 329654 0 329710 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 332690 0 332746 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 335726 0 335782 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 338762 0 338818 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 147494 0 147550 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 341798 0 341854 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 344834 0 344890 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 347870 0 347926 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 350906 0 350962 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 353942 0 353998 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 356978 0 357034 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 360014 0 360070 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 363050 0 363106 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 366086 0 366142 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 369122 0 369178 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 150530 0 150586 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 372158 0 372214 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 375194 0 375250 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 378230 0 378286 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 381266 0 381322 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 384302 0 384358 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 387338 0 387394 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 390374 0 390430 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 393410 0 393466 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 396446 0 396502 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 399482 0 399538 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 153566 0 153622 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 402518 0 402574 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 405554 0 405610 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 408590 0 408646 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 411626 0 411682 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 414662 0 414718 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 417698 0 417754 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 420734 0 420790 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 423770 0 423826 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 426806 0 426862 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 429842 0 429898 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 156602 0 156658 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 130290 0 130346 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 433890 0 433946 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 436926 0 436982 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 439962 0 440018 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 442998 0 443054 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 446034 0 446090 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 449070 0 449126 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 452106 0 452162 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 455142 0 455198 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 458178 0 458234 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 461214 0 461270 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 160650 0 160706 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 464250 0 464306 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 467286 0 467342 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 470322 0 470378 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 473358 0 473414 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 476394 0 476450 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 479430 0 479486 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 482466 0 482522 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 485502 0 485558 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 488538 0 488594 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 491574 0 491630 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 163686 0 163742 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 494610 0 494666 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 497646 0 497702 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 500682 0 500738 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 503718 0 503774 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 506754 0 506810 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 509790 0 509846 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 512826 0 512882 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 515862 0 515918 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 166722 0 166778 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 169758 0 169814 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 172794 0 172850 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 175830 0 175886 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 178866 0 178922 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 181902 0 181958 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 184938 0 184994 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 187974 0 188030 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 133326 0 133382 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 191010 0 191066 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 194046 0 194102 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 197082 0 197138 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 200118 0 200174 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 203154 0 203210 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 206190 0 206246 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 209226 0 209282 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 212262 0 212318 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 215298 0 215354 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 218334 0 218390 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 136362 0 136418 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 221370 0 221426 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 224406 0 224462 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 227442 0 227498 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 230478 0 230534 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 233514 0 233570 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 236550 0 236606 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 239586 0 239642 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 242622 0 242678 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 245658 0 245714 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 248694 0 248750 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 139398 0 139454 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 251730 0 251786 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 254766 0 254822 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 257802 0 257858 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 260838 0 260894 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 263874 0 263930 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 266910 0 266966 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 269946 0 270002 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 272982 0 273038 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 276018 0 276074 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 279054 0 279110 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 142434 0 142490 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 282090 0 282146 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 285126 0 285182 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 288162 0 288218 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 291198 0 291254 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 294234 0 294290 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 297270 0 297326 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 300306 0 300362 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 303342 0 303398 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 306378 0 306434 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 309414 0 309470 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 145470 0 145526 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 312450 0 312506 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 315486 0 315542 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 318522 0 318578 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 321558 0 321614 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 324594 0 324650 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 327630 0 327686 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 330666 0 330722 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 333702 0 333758 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 336738 0 336794 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 339774 0 339830 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 148506 0 148562 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 342810 0 342866 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 345846 0 345902 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 348882 0 348938 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 351918 0 351974 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 354954 0 355010 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 357990 0 358046 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 361026 0 361082 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 364062 0 364118 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 367098 0 367154 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 370134 0 370190 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 151542 0 151598 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 373170 0 373226 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 376206 0 376262 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 379242 0 379298 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 382278 0 382334 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 385314 0 385370 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 388350 0 388406 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 391386 0 391442 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 394422 0 394478 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 397458 0 397514 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 400494 0 400550 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 154578 0 154634 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 403530 0 403586 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 406566 0 406622 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 409602 0 409658 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 412638 0 412694 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 415674 0 415730 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 418710 0 418766 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 421746 0 421802 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 424782 0 424838 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 427818 0 427874 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 430854 0 430910 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 157614 0 157670 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 317744 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 317744 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 317744 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 317744 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 317744 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 317744 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 317744 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 317744 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 317744 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 317744 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 317744 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 317744 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 372848 2128 373168 317744 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 403568 2128 403888 317744 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 434288 2128 434608 317744 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 465008 2128 465328 317744 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 495728 2128 496048 317744 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 526448 2128 526768 317744 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 317744 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 317744 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 317744 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 317744 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 317744 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 317744 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 317744 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 317744 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 317744 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 317744 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 317744 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 357488 2128 357808 317744 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 388208 2128 388528 317744 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 418928 2128 419248 317744 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 449648 2128 449968 317744 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 480368 2128 480688 317744 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 511088 2128 511408 317744 6 vssd1
port 503 nsew ground bidirectional
rlabel metal2 s 20994 0 21050 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 22006 0 22062 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 23018 0 23074 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 27066 0 27122 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 61474 0 61530 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 64510 0 64566 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 67546 0 67602 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 70582 0 70638 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 73618 0 73674 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 76654 0 76710 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 79690 0 79746 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 82726 0 82782 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 85762 0 85818 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 88798 0 88854 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 31114 0 31170 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 91834 0 91890 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 94870 0 94926 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 97906 0 97962 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 100942 0 100998 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 103978 0 104034 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 107014 0 107070 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 110050 0 110106 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 113086 0 113142 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 116122 0 116178 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 119158 0 119214 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 35162 0 35218 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 122194 0 122250 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 125230 0 125286 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 39210 0 39266 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 43258 0 43314 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 46294 0 46350 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 49330 0 49386 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 52366 0 52422 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 58438 0 58494 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 24030 0 24086 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 62486 0 62542 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 65522 0 65578 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 68558 0 68614 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 71594 0 71650 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 74630 0 74686 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 77666 0 77722 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 80702 0 80758 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 83738 0 83794 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 86774 0 86830 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 89810 0 89866 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 32126 0 32182 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 92846 0 92902 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 95882 0 95938 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 98918 0 98974 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 101954 0 102010 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 104990 0 105046 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 108026 0 108082 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 111062 0 111118 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 114098 0 114154 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 117134 0 117190 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 120170 0 120226 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 36174 0 36230 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 123206 0 123262 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 126242 0 126298 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 40222 0 40278 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 44270 0 44326 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 47306 0 47362 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 50342 0 50398 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 53378 0 53434 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 56414 0 56470 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 59450 0 59506 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 29090 0 29146 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 63498 0 63554 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 66534 0 66590 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 69570 0 69626 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 72606 0 72662 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 75642 0 75698 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 78678 0 78734 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 81714 0 81770 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 84750 0 84806 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 87786 0 87842 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 90822 0 90878 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 33138 0 33194 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 93858 0 93914 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 96894 0 96950 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 99930 0 99986 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 102966 0 103022 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 106002 0 106058 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 109038 0 109094 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 112074 0 112130 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 115110 0 115166 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 118146 0 118202 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 121182 0 121238 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 37186 0 37242 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 124218 0 124274 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 127254 0 127310 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 41234 0 41290 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 45282 0 45338 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 48318 0 48374 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 51354 0 51410 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 54390 0 54446 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 57426 0 57482 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 60462 0 60518 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 30102 0 30158 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 38198 0 38254 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 42246 0 42302 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 25042 0 25098 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 26054 0 26110 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 540000 320000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 86939898
string GDS_FILE /home/anton/projects/CUP-algofoogle/openlane/user_proj_example/runs/24_09_24_09_37/results/signoff/user_proj_example.magic.gds
string GDS_START 1381882
<< end >>

